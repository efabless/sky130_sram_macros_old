VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_8kbyte_1rw1r_32x2048_8
   CLASS BLOCK ;
   SIZE 1080.22 BY 709.62 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.96 0.0 117.34 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  123.76 0.0 124.14 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  129.2 0.0 129.58 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  135.32 0.0 135.7 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  140.08 0.0 140.46 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  146.88 0.0 147.26 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  152.32 0.0 152.7 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.76 0.0 158.14 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.88 0.0 164.26 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  169.32 0.0 169.7 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  176.12 0.0 176.5 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  181.56 0.0 181.94 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  187.0 0.0 187.38 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  193.12 0.0 193.5 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  198.56 0.0 198.94 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 0.0 205.74 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  210.8 0.0 211.18 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  216.92 0.0 217.3 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  223.04 0.0 223.42 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  228.48 0.0 228.86 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  233.92 0.0 234.3 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  239.36 0.0 239.74 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  245.48 0.0 245.86 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  251.6 0.0 251.98 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  257.72 0.0 258.1 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  263.16 0.0 263.54 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  268.6 0.0 268.98 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.72 0.0 275.1 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  280.84 0.0 281.22 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  286.96 0.0 287.34 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  293.08 0.0 293.46 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 0.0 298.22 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  76.16 0.0 76.54 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  82.28 0.0 82.66 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.72 0.0 88.1 0.38 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 168.64 0.38 169.02 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 176.8 0.38 177.18 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 183.6 0.38 183.98 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 191.76 0.38 192.14 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 197.2 0.38 197.58 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 205.36 0.38 205.74 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 210.8 0.38 211.18 ;
      END
   END addr0[9]
   PIN addr0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 220.32 0.38 220.7 ;
      END
   END addr0[10]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  998.92 709.24 999.3 709.62 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  993.48 709.24 993.86 709.62 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  986.68 709.24 987.06 709.62 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1079.84 115.6 1080.22 115.98 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1079.84 107.44 1080.22 107.82 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1079.84 102.0 1080.22 102.38 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1079.84 92.48 1080.22 92.86 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1079.84 87.04 1080.22 87.42 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1079.84 78.88 1080.22 79.26 ;
      END
   END addr1[8]
   PIN addr1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1079.84 72.76 1080.22 73.14 ;
      END
   END addr1[9]
   PIN addr1[10]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1079.84 64.6 1080.22 64.98 ;
      END
   END addr1[10]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 59.84 0.38 60.22 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1079.84 668.44 1080.22 668.82 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 68.68 0.38 69.06 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 61.2 0.38 61.58 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1079.84 667.08 1080.22 667.46 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.84 0.0 94.22 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  99.28 0.0 99.66 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  105.4 0.0 105.78 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  111.52 0.0 111.9 0.38 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  138.72 0.0 139.1 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.6 0.0 166.98 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.08 0.0 191.46 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  214.88 0.0 215.26 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 0.0 241.78 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  266.56 0.0 266.94 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  290.36 0.0 290.74 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.2 0.0 316.58 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  341.36 0.0 341.74 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  365.84 0.0 366.22 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  391.0 0.0 391.38 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  415.48 0.0 415.86 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  440.64 0.0 441.02 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  465.8 0.0 466.18 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  490.96 0.0 491.34 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  515.44 0.0 515.82 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  539.24 0.0 539.62 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  565.76 0.0 566.14 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  590.24 0.0 590.62 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  615.4 0.0 615.78 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  640.56 0.0 640.94 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  665.72 0.0 666.1 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  690.2 0.0 690.58 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  715.36 0.0 715.74 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  739.16 0.0 739.54 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  765.0 0.0 765.38 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  790.16 0.0 790.54 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  815.32 0.0 815.7 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  839.8 0.0 840.18 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  864.96 0.0 865.34 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  890.12 0.0 890.5 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  915.28 0.0 915.66 0.38 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  141.44 709.24 141.82 709.62 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  165.92 709.24 166.3 709.62 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.08 709.24 191.46 709.62 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.24 709.24 216.62 709.62 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 709.24 241.78 709.62 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  266.56 709.24 266.94 709.62 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  291.04 709.24 291.42 709.62 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.2 709.24 316.58 709.62 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  341.36 709.24 341.74 709.62 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  366.52 709.24 366.9 709.62 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  391.68 709.24 392.06 709.62 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  415.48 709.24 415.86 709.62 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  440.64 709.24 441.02 709.62 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  466.48 709.24 466.86 709.62 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  490.96 709.24 491.34 709.62 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  515.44 709.24 515.82 709.62 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  540.6 709.24 540.98 709.62 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  565.76 709.24 566.14 709.62 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  590.24 709.24 590.62 709.62 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  615.4 709.24 615.78 709.62 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  640.56 709.24 640.94 709.62 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  665.72 709.24 666.1 709.62 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  690.88 709.24 691.26 709.62 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  715.36 709.24 715.74 709.62 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  740.52 709.24 740.9 709.62 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  765.68 709.24 766.06 709.62 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  790.84 709.24 791.22 709.62 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  816.0 709.24 816.38 709.62 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  839.8 709.24 840.18 709.62 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  864.96 709.24 865.34 709.62 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  890.8 709.24 891.18 709.62 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  915.28 709.24 915.66 709.62 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  1.36 0.0 2.42 708.94 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.06 708.94 ;
      END
   END gnd
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 1079.6 709.0 ;
   LAYER  met2 ;
      RECT  0.62 0.62 1079.6 709.0 ;
   LAYER  met3 ;
      RECT  0.68 168.34 1079.6 169.32 ;
      RECT  0.62 169.32 0.68 176.5 ;
      RECT  0.62 177.48 0.68 183.3 ;
      RECT  0.62 184.28 0.68 191.46 ;
      RECT  0.62 192.44 0.68 196.9 ;
      RECT  0.62 197.88 0.68 205.06 ;
      RECT  0.62 206.04 0.68 210.5 ;
      RECT  0.62 211.48 0.68 220.02 ;
      RECT  0.62 221.0 0.68 709.0 ;
      RECT  0.68 0.62 1079.54 115.3 ;
      RECT  0.68 115.3 1079.54 116.28 ;
      RECT  0.68 116.28 1079.54 168.34 ;
      RECT  1079.54 116.28 1079.6 168.34 ;
      RECT  1079.54 108.12 1079.6 115.3 ;
      RECT  1079.54 102.68 1079.6 107.14 ;
      RECT  1079.54 93.16 1079.6 101.7 ;
      RECT  1079.54 87.72 1079.6 92.18 ;
      RECT  1079.54 79.56 1079.6 86.74 ;
      RECT  1079.54 73.44 1079.6 78.58 ;
      RECT  1079.54 0.62 1079.6 64.3 ;
      RECT  1079.54 65.28 1079.6 72.46 ;
      RECT  0.62 0.62 0.68 59.54 ;
      RECT  0.68 169.32 1079.54 668.14 ;
      RECT  0.68 668.14 1079.54 669.12 ;
      RECT  0.68 669.12 1079.54 709.0 ;
      RECT  1079.54 669.12 1079.6 709.0 ;
      RECT  0.62 69.36 0.68 168.34 ;
      RECT  0.62 60.52 0.68 60.9 ;
      RECT  0.62 61.88 0.68 68.38 ;
      RECT  1079.54 169.32 1079.6 666.78 ;
      RECT  1079.54 667.76 1079.6 668.14 ;
   LAYER  met4 ;
      RECT  116.66 0.68 117.64 709.0 ;
      RECT  117.64 0.62 123.46 0.68 ;
      RECT  124.44 0.62 128.9 0.68 ;
      RECT  129.88 0.62 135.02 0.68 ;
      RECT  140.76 0.62 146.58 0.68 ;
      RECT  147.56 0.62 152.02 0.68 ;
      RECT  153.0 0.62 157.46 0.68 ;
      RECT  158.44 0.62 163.58 0.68 ;
      RECT  170.0 0.62 175.82 0.68 ;
      RECT  176.8 0.62 181.26 0.68 ;
      RECT  182.24 0.62 186.7 0.68 ;
      RECT  193.8 0.62 198.26 0.68 ;
      RECT  199.24 0.62 205.06 0.68 ;
      RECT  206.04 0.62 210.5 0.68 ;
      RECT  217.6 0.62 222.74 0.68 ;
      RECT  223.72 0.62 228.18 0.68 ;
      RECT  229.16 0.62 233.62 0.68 ;
      RECT  234.6 0.62 239.06 0.68 ;
      RECT  246.16 0.62 251.3 0.68 ;
      RECT  252.28 0.62 257.42 0.68 ;
      RECT  258.4 0.62 262.86 0.68 ;
      RECT  269.28 0.62 274.42 0.68 ;
      RECT  275.4 0.62 280.54 0.68 ;
      RECT  281.52 0.62 286.66 0.68 ;
      RECT  293.76 0.62 297.54 0.68 ;
      RECT  76.84 0.62 81.98 0.68 ;
      RECT  82.96 0.62 87.42 0.68 ;
      RECT  117.64 0.68 998.62 708.94 ;
      RECT  998.62 0.68 999.6 708.94 ;
      RECT  999.6 0.68 1079.6 708.94 ;
      RECT  999.6 708.94 1079.6 709.0 ;
      RECT  994.16 708.94 998.62 709.0 ;
      RECT  987.36 708.94 993.18 709.0 ;
      RECT  88.4 0.62 93.54 0.68 ;
      RECT  94.52 0.62 98.98 0.68 ;
      RECT  99.96 0.62 105.1 0.68 ;
      RECT  106.08 0.62 111.22 0.68 ;
      RECT  112.2 0.62 116.66 0.68 ;
      RECT  136.0 0.62 138.42 0.68 ;
      RECT  139.4 0.62 139.78 0.68 ;
      RECT  164.56 0.62 166.3 0.68 ;
      RECT  167.28 0.62 169.02 0.68 ;
      RECT  187.68 0.62 190.78 0.68 ;
      RECT  191.76 0.62 192.82 0.68 ;
      RECT  211.48 0.62 214.58 0.68 ;
      RECT  215.56 0.62 216.62 0.68 ;
      RECT  240.04 0.62 241.1 0.68 ;
      RECT  242.08 0.62 245.18 0.68 ;
      RECT  263.84 0.62 266.26 0.68 ;
      RECT  267.24 0.62 268.3 0.68 ;
      RECT  287.64 0.62 290.06 0.68 ;
      RECT  291.04 0.62 292.78 0.68 ;
      RECT  298.52 0.62 315.9 0.68 ;
      RECT  316.88 0.62 341.06 0.68 ;
      RECT  342.04 0.62 365.54 0.68 ;
      RECT  366.52 0.62 390.7 0.68 ;
      RECT  391.68 0.62 415.18 0.68 ;
      RECT  416.16 0.62 440.34 0.68 ;
      RECT  441.32 0.62 465.5 0.68 ;
      RECT  466.48 0.62 490.66 0.68 ;
      RECT  491.64 0.62 515.14 0.68 ;
      RECT  516.12 0.62 538.94 0.68 ;
      RECT  539.92 0.62 565.46 0.68 ;
      RECT  566.44 0.62 589.94 0.68 ;
      RECT  590.92 0.62 615.1 0.68 ;
      RECT  616.08 0.62 640.26 0.68 ;
      RECT  641.24 0.62 665.42 0.68 ;
      RECT  666.4 0.62 689.9 0.68 ;
      RECT  690.88 0.62 715.06 0.68 ;
      RECT  716.04 0.62 738.86 0.68 ;
      RECT  739.84 0.62 764.7 0.68 ;
      RECT  765.68 0.62 789.86 0.68 ;
      RECT  790.84 0.62 815.02 0.68 ;
      RECT  816.0 0.62 839.5 0.68 ;
      RECT  840.48 0.62 864.66 0.68 ;
      RECT  865.64 0.62 889.82 0.68 ;
      RECT  890.8 0.62 914.98 0.68 ;
      RECT  915.96 0.62 1079.6 0.68 ;
      RECT  117.64 708.94 141.14 709.0 ;
      RECT  142.12 708.94 165.62 709.0 ;
      RECT  166.6 708.94 190.78 709.0 ;
      RECT  191.76 708.94 215.94 709.0 ;
      RECT  216.92 708.94 241.1 709.0 ;
      RECT  242.08 708.94 266.26 709.0 ;
      RECT  267.24 708.94 290.74 709.0 ;
      RECT  291.72 708.94 315.9 709.0 ;
      RECT  316.88 708.94 341.06 709.0 ;
      RECT  342.04 708.94 366.22 709.0 ;
      RECT  367.2 708.94 391.38 709.0 ;
      RECT  392.36 708.94 415.18 709.0 ;
      RECT  416.16 708.94 440.34 709.0 ;
      RECT  441.32 708.94 466.18 709.0 ;
      RECT  467.16 708.94 490.66 709.0 ;
      RECT  491.64 708.94 515.14 709.0 ;
      RECT  516.12 708.94 540.3 709.0 ;
      RECT  541.28 708.94 565.46 709.0 ;
      RECT  566.44 708.94 589.94 709.0 ;
      RECT  590.92 708.94 615.1 709.0 ;
      RECT  616.08 708.94 640.26 709.0 ;
      RECT  641.24 708.94 665.42 709.0 ;
      RECT  666.4 708.94 690.58 709.0 ;
      RECT  691.56 708.94 715.06 709.0 ;
      RECT  716.04 708.94 740.22 709.0 ;
      RECT  741.2 708.94 765.38 709.0 ;
      RECT  766.36 708.94 790.54 709.0 ;
      RECT  791.52 708.94 815.7 709.0 ;
      RECT  816.68 708.94 839.5 709.0 ;
      RECT  840.48 708.94 864.66 709.0 ;
      RECT  865.64 708.94 890.5 709.0 ;
      RECT  891.48 708.94 914.98 709.0 ;
      RECT  915.96 708.94 986.38 709.0 ;
      RECT  2.72 0.68 116.66 709.0 ;
      RECT  2.72 0.62 75.86 0.68 ;
   END
END    sky130_sram_8kbyte_1rw1r_32x2048_8
END    LIBRARY
