VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_4kbyte_1rw1r_32x1024_8
   CLASS BLOCK ;
   SIZE 670.86 BY 651.14 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  106.76 0.0 107.14 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  112.2 0.0 112.58 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  118.32 0.0 118.7 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  123.76 0.0 124.14 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  129.2 0.0 129.58 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  134.64 0.0 135.02 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  141.44 0.0 141.82 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  147.56 0.0 147.94 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  153.0 0.0 153.38 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  158.44 0.0 158.82 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.88 0.0 164.26 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  170.68 0.0 171.06 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  176.12 0.0 176.5 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  181.56 0.0 181.94 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  188.36 0.0 188.74 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  194.48 0.0 194.86 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  199.92 0.0 200.3 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 0.0 205.74 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  210.8 0.0 211.18 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 0.0 217.98 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  223.04 0.0 223.42 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  229.16 0.0 229.54 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  234.6 0.0 234.98 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  240.04 0.0 240.42 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  246.84 0.0 247.22 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  252.28 0.0 252.66 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  257.72 0.0 258.1 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  263.16 0.0 263.54 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  269.96 0.0 270.34 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 0.0 276.46 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  281.52 0.0 281.9 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  286.96 0.0 287.34 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  71.4 0.0 71.78 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  76.84 0.0 77.22 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 140.08 0.38 140.46 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 148.24 0.38 148.62 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 155.04 0.38 155.42 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 162.52 0.38 162.9 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 167.96 0.38 168.34 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 176.8 0.38 177.18 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 182.24 0.38 182.62 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 191.76 0.38 192.14 ;
      END
   END addr0[9]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  594.32 650.76 594.7 651.14 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  588.2 650.76 588.58 651.14 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  670.48 83.64 670.86 84.02 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  670.48 75.48 670.86 75.86 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  670.48 69.36 670.86 69.74 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  670.48 61.2 670.86 61.58 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  610.64 0.0 611.02 0.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  612.68 0.0 613.06 0.38 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  611.32 0.0 611.7 0.38 ;
      END
   END addr1[8]
   PIN addr1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  612.0 0.0 612.38 0.38 ;
      END
   END addr1[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 31.28 0.38 31.66 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  670.48 639.88 670.86 640.26 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 40.8 0.38 41.18 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 32.64 0.38 33.02 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  652.12 650.76 652.5 651.14 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  82.28 0.0 82.66 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  89.08 0.0 89.46 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.84 0.0 94.22 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  99.96 0.0 100.34 0.38 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  133.28 0.0 133.66 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.24 0.0 148.62 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.48 0.0 160.86 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.4 0.0 173.78 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  185.64 0.0 186.02 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 0.0 197.58 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.44 0.0 209.82 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  221.0 0.0 221.38 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  238.0 0.0 238.38 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.2 0.0 248.58 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  261.12 0.0 261.5 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  273.36 0.0 273.74 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 0.0 285.3 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 0.0 298.22 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  310.76 0.0 311.14 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  323.0 0.0 323.38 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  335.92 0.0 336.3 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  348.16 0.0 348.54 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  360.4 0.0 360.78 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  372.64 0.0 373.02 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  385.56 0.0 385.94 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  397.8 0.0 398.18 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  410.04 0.0 410.42 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  422.96 0.0 423.34 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  433.84 0.0 434.22 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  448.12 0.0 448.5 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  460.36 0.0 460.74 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  472.6 0.0 472.98 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  485.52 0.0 485.9 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  497.76 0.0 498.14 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  510.0 0.0 510.38 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  522.92 0.0 523.3 0.38 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  136.68 650.76 137.06 651.14 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.24 650.76 148.62 651.14 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  161.16 650.76 161.54 651.14 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.4 650.76 173.78 651.14 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.32 650.76 186.7 651.14 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.56 650.76 198.94 651.14 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  211.48 650.76 211.86 651.14 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.72 650.76 224.1 651.14 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.96 650.76 236.34 651.14 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.2 650.76 248.58 651.14 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  260.44 650.76 260.82 651.14 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  273.36 650.76 273.74 651.14 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  286.28 650.76 286.66 651.14 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  298.52 650.76 298.9 651.14 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  311.44 650.76 311.82 651.14 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  323.68 650.76 324.06 651.14 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  335.24 650.76 335.62 651.14 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  348.84 650.76 349.22 651.14 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  360.4 650.76 360.78 651.14 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  373.32 650.76 373.7 651.14 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  385.56 650.76 385.94 651.14 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  398.48 650.76 398.86 651.14 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  410.72 650.76 411.1 651.14 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  423.64 650.76 424.02 651.14 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  435.88 650.76 436.26 651.14 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  448.12 650.76 448.5 651.14 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  460.36 650.76 460.74 651.14 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  472.6 650.76 472.98 651.14 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  485.52 650.76 485.9 651.14 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  498.44 650.76 498.82 651.14 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  510.68 650.76 511.06 651.14 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  523.6 650.76 523.98 651.14 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 35.36 0.6 36.42 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 28.56 0.6 29.62 ;
      END
   END gnd
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 670.24 650.52 ;
   LAYER  met2 ;
      RECT  0.62 0.62 670.24 650.52 ;
   LAYER  met3 ;
      RECT  0.68 139.78 670.24 140.76 ;
      RECT  0.62 140.76 0.68 147.94 ;
      RECT  0.62 148.92 0.68 154.74 ;
      RECT  0.62 155.72 0.68 162.22 ;
      RECT  0.62 163.2 0.68 167.66 ;
      RECT  0.62 168.64 0.68 176.5 ;
      RECT  0.62 177.48 0.68 181.94 ;
      RECT  0.62 182.92 0.68 191.46 ;
      RECT  0.62 192.44 0.68 650.52 ;
      RECT  0.68 83.34 670.18 84.32 ;
      RECT  0.68 84.32 670.18 139.78 ;
      RECT  670.18 84.32 670.24 139.78 ;
      RECT  670.18 76.16 670.24 83.34 ;
      RECT  670.18 70.04 670.24 75.18 ;
      RECT  670.18 0.62 670.24 60.9 ;
      RECT  670.18 61.88 670.24 69.06 ;
      RECT  0.68 140.76 670.18 639.58 ;
      RECT  0.68 639.58 670.18 640.56 ;
      RECT  0.68 640.56 670.18 650.52 ;
      RECT  670.18 140.76 670.24 639.58 ;
      RECT  670.18 640.56 670.24 650.52 ;
      RECT  0.62 41.48 0.68 139.78 ;
      RECT  0.62 31.96 0.68 32.34 ;
      RECT  0.68 36.72 0.9 83.34 ;
      RECT  0.9 0.62 670.18 35.06 ;
      RECT  0.9 35.06 670.18 36.72 ;
      RECT  0.9 36.72 670.18 83.34 ;
      RECT  0.62 33.32 0.68 35.06 ;
      RECT  0.62 36.72 0.68 40.5 ;
      RECT  0.62 0.62 0.68 28.26 ;
      RECT  0.62 29.92 0.68 30.98 ;
      RECT  0.68 0.62 0.9 28.26 ;
      RECT  0.68 29.92 0.9 35.06 ;
   LAYER  met4 ;
      RECT  0.62 0.68 106.46 650.52 ;
      RECT  106.46 0.68 107.44 650.52 ;
      RECT  107.44 0.62 111.9 0.68 ;
      RECT  112.88 0.62 118.02 0.68 ;
      RECT  119.0 0.62 123.46 0.68 ;
      RECT  124.44 0.62 128.9 0.68 ;
      RECT  135.32 0.62 141.14 0.68 ;
      RECT  142.12 0.62 147.26 0.68 ;
      RECT  153.68 0.62 158.14 0.68 ;
      RECT  164.56 0.62 170.38 0.68 ;
      RECT  176.8 0.62 181.26 0.68 ;
      RECT  189.04 0.62 194.18 0.68 ;
      RECT  200.6 0.62 205.06 0.68 ;
      RECT  211.48 0.62 217.3 0.68 ;
      RECT  223.72 0.62 228.86 0.68 ;
      RECT  229.84 0.62 234.3 0.68 ;
      RECT  240.72 0.62 246.54 0.68 ;
      RECT  252.96 0.62 257.42 0.68 ;
      RECT  263.84 0.62 269.66 0.68 ;
      RECT  276.76 0.62 281.22 0.68 ;
      RECT  0.62 0.62 71.1 0.68 ;
      RECT  72.08 0.62 76.54 0.68 ;
      RECT  107.44 0.68 594.02 650.46 ;
      RECT  594.02 0.68 595.0 650.46 ;
      RECT  595.0 0.68 670.24 650.46 ;
      RECT  588.88 650.46 594.02 650.52 ;
      RECT  613.36 0.62 670.24 0.68 ;
      RECT  595.0 650.46 651.82 650.52 ;
      RECT  652.8 650.46 670.24 650.52 ;
      RECT  77.52 0.62 81.98 0.68 ;
      RECT  82.96 0.62 88.78 0.68 ;
      RECT  89.76 0.62 93.54 0.68 ;
      RECT  94.52 0.62 99.66 0.68 ;
      RECT  100.64 0.62 106.46 0.68 ;
      RECT  129.88 0.62 132.98 0.68 ;
      RECT  133.96 0.62 134.34 0.68 ;
      RECT  148.92 0.62 152.7 0.68 ;
      RECT  159.12 0.62 160.18 0.68 ;
      RECT  161.16 0.62 163.58 0.68 ;
      RECT  171.36 0.62 173.1 0.68 ;
      RECT  174.08 0.62 175.82 0.68 ;
      RECT  182.24 0.62 185.34 0.68 ;
      RECT  186.32 0.62 188.06 0.68 ;
      RECT  195.16 0.62 196.9 0.68 ;
      RECT  197.88 0.62 199.62 0.68 ;
      RECT  206.04 0.62 209.14 0.68 ;
      RECT  210.12 0.62 210.5 0.68 ;
      RECT  218.28 0.62 220.7 0.68 ;
      RECT  221.68 0.62 222.74 0.68 ;
      RECT  235.28 0.62 237.7 0.68 ;
      RECT  238.68 0.62 239.74 0.68 ;
      RECT  247.52 0.62 247.9 0.68 ;
      RECT  248.88 0.62 251.98 0.68 ;
      RECT  258.4 0.62 260.82 0.68 ;
      RECT  261.8 0.62 262.86 0.68 ;
      RECT  270.64 0.62 273.06 0.68 ;
      RECT  274.04 0.62 275.78 0.68 ;
      RECT  282.2 0.62 284.62 0.68 ;
      RECT  285.6 0.62 286.66 0.68 ;
      RECT  287.64 0.62 297.54 0.68 ;
      RECT  298.52 0.62 310.46 0.68 ;
      RECT  311.44 0.62 322.7 0.68 ;
      RECT  323.68 0.62 335.62 0.68 ;
      RECT  336.6 0.62 347.86 0.68 ;
      RECT  348.84 0.62 360.1 0.68 ;
      RECT  361.08 0.62 372.34 0.68 ;
      RECT  373.32 0.62 385.26 0.68 ;
      RECT  386.24 0.62 397.5 0.68 ;
      RECT  398.48 0.62 409.74 0.68 ;
      RECT  410.72 0.62 422.66 0.68 ;
      RECT  423.64 0.62 433.54 0.68 ;
      RECT  434.52 0.62 447.82 0.68 ;
      RECT  448.8 0.62 460.06 0.68 ;
      RECT  461.04 0.62 472.3 0.68 ;
      RECT  473.28 0.62 485.22 0.68 ;
      RECT  486.2 0.62 497.46 0.68 ;
      RECT  498.44 0.62 509.7 0.68 ;
      RECT  510.68 0.62 522.62 0.68 ;
      RECT  523.6 0.62 610.34 0.68 ;
      RECT  107.44 650.46 136.38 650.52 ;
      RECT  137.36 650.46 147.94 650.52 ;
      RECT  148.92 650.46 160.86 650.52 ;
      RECT  161.84 650.46 173.1 650.52 ;
      RECT  174.08 650.46 186.02 650.52 ;
      RECT  187.0 650.46 198.26 650.52 ;
      RECT  199.24 650.46 211.18 650.52 ;
      RECT  212.16 650.46 223.42 650.52 ;
      RECT  224.4 650.46 235.66 650.52 ;
      RECT  236.64 650.46 247.9 650.52 ;
      RECT  248.88 650.46 260.14 650.52 ;
      RECT  261.12 650.46 273.06 650.52 ;
      RECT  274.04 650.46 285.98 650.52 ;
      RECT  286.96 650.46 298.22 650.52 ;
      RECT  299.2 650.46 311.14 650.52 ;
      RECT  312.12 650.46 323.38 650.52 ;
      RECT  324.36 650.46 334.94 650.52 ;
      RECT  335.92 650.46 348.54 650.52 ;
      RECT  349.52 650.46 360.1 650.52 ;
      RECT  361.08 650.46 373.02 650.52 ;
      RECT  374.0 650.46 385.26 650.52 ;
      RECT  386.24 650.46 398.18 650.52 ;
      RECT  399.16 650.46 410.42 650.52 ;
      RECT  411.4 650.46 423.34 650.52 ;
      RECT  424.32 650.46 435.58 650.52 ;
      RECT  436.56 650.46 447.82 650.52 ;
      RECT  448.8 650.46 460.06 650.52 ;
      RECT  461.04 650.46 472.3 650.52 ;
      RECT  473.28 650.46 485.22 650.52 ;
      RECT  486.2 650.46 498.14 650.52 ;
      RECT  499.12 650.46 510.38 650.52 ;
      RECT  511.36 650.46 523.3 650.52 ;
      RECT  524.28 650.46 587.9 650.52 ;
   END
END    sky130_sram_4kbyte_1rw1r_32x1024_8
END    LIBRARY
