VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_1kbyte_1rw1r_8x1024_8
   CLASS BLOCK ;
   SIZE 451.9 BY 443.06 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.04 0.0 87.42 0.64 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.16 0.0 93.54 0.64 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  98.6 0.0 98.98 0.64 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.04 0.0 104.42 0.64 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.16 0.0 110.54 0.64 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  115.6 0.0 115.98 0.64 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  122.4 0.0 122.78 0.64 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.16 0.0 127.54 0.64 ;
      END
   END din0[7]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  63.24 0.0 63.62 0.64 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  70.04 0.0 70.42 0.64 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  75.48 0.0 75.86 0.64 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 141.44 0.64 141.82 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 149.6 0.64 149.98 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 156.4 0.64 156.78 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 164.56 0.64 164.94 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 169.32 0.64 169.7 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 177.48 0.64 177.86 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 183.6 0.64 183.98 ;
      END
   END addr0[9]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  382.16 442.42 382.54 443.06 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  376.72 442.42 377.1 443.06 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  371.28 442.42 371.66 443.06 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  451.26 97.24 451.9 97.62 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  451.26 88.4 451.9 88.78 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  451.26 82.96 451.9 83.34 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  451.26 74.12 451.9 74.5 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  451.26 68.68 451.9 69.06 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  451.26 59.84 451.9 60.22 ;
      END
   END addr1[8]
   PIN addr1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  451.26 53.72 451.9 54.1 ;
      END
   END addr1[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 41.48 0.64 41.86 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  451.26 395.76 451.9 396.14 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 49.64 0.64 50.02 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 42.16 0.64 42.54 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  451.26 395.08 451.9 395.46 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.92 0.0 81.3 0.64 ;
      END
   END wmask0[0]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  125.12 0.0 125.5 0.64 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  150.96 0.0 151.34 0.64 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.12 0.0 176.5 0.64 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.28 0.0 201.66 0.64 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  226.44 0.0 226.82 0.64 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 0.0 251.3 0.64 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 0.0 276.46 0.64 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  301.24 0.0 301.62 0.64 ;
      END
   END dout0[7]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  126.48 442.42 126.86 443.06 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  151.64 442.42 152.02 443.06 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.8 442.42 177.18 443.06 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.96 442.42 202.34 443.06 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  226.44 442.42 226.82 443.06 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 442.42 251.3 443.06 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.76 442.42 277.14 443.06 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  301.92 442.42 302.3 443.06 ;
      END
   END dout1[7]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  448.8 1.36 450.54 441.7 ;
         LAYER met3 ;
         RECT  1.36 439.96 450.54 441.7 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 441.7 ;
         LAYER met3 ;
         RECT  1.36 1.36 450.54 3.1 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  4.76 4.76 447.14 6.5 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 438.3 ;
         LAYER met3 ;
         RECT  4.76 436.56 447.14 438.3 ;
         LAYER met4 ;
         RECT  445.4 4.76 447.14 438.3 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 451.28 442.44 ;
   LAYER  met2 ;
      RECT  0.62 0.62 451.28 442.44 ;
   LAYER  met3 ;
      RECT  0.98 140.84 451.28 142.42 ;
      RECT  0.62 142.42 0.98 149.0 ;
      RECT  0.62 150.58 0.98 155.8 ;
      RECT  0.62 157.38 0.98 163.96 ;
      RECT  0.62 165.54 0.98 168.72 ;
      RECT  0.62 170.3 0.98 176.88 ;
      RECT  0.62 178.46 0.98 183.0 ;
      RECT  0.98 96.64 450.92 98.22 ;
      RECT  0.98 98.22 450.92 140.84 ;
      RECT  450.92 98.22 451.28 140.84 ;
      RECT  450.92 89.38 451.28 96.64 ;
      RECT  450.92 83.94 451.28 87.8 ;
      RECT  450.92 75.1 451.28 82.36 ;
      RECT  450.92 69.66 451.28 73.52 ;
      RECT  450.92 60.82 451.28 68.08 ;
      RECT  450.92 54.7 451.28 59.24 ;
      RECT  0.98 142.42 450.92 395.16 ;
      RECT  0.98 395.16 450.92 396.74 ;
      RECT  0.62 50.62 0.98 140.84 ;
      RECT  0.62 43.14 0.98 49.04 ;
      RECT  450.92 142.42 451.28 394.48 ;
      RECT  0.62 184.58 0.76 439.36 ;
      RECT  0.62 439.36 0.76 442.3 ;
      RECT  0.62 442.3 0.76 442.44 ;
      RECT  0.76 184.58 0.98 439.36 ;
      RECT  0.76 442.3 0.98 442.44 ;
      RECT  0.98 442.3 450.92 442.44 ;
      RECT  450.92 396.74 451.14 439.36 ;
      RECT  450.92 442.3 451.14 442.44 ;
      RECT  451.14 396.74 451.28 439.36 ;
      RECT  451.14 439.36 451.28 442.3 ;
      RECT  451.14 442.3 451.28 442.44 ;
      RECT  0.98 0.62 450.92 0.76 ;
      RECT  450.92 0.62 451.14 0.76 ;
      RECT  450.92 3.7 451.14 53.12 ;
      RECT  451.14 0.62 451.28 0.76 ;
      RECT  451.14 0.76 451.28 3.7 ;
      RECT  451.14 3.7 451.28 53.12 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 40.88 ;
      RECT  0.76 0.62 0.98 0.76 ;
      RECT  0.76 3.7 0.98 40.88 ;
      RECT  0.98 3.7 4.16 4.16 ;
      RECT  0.98 4.16 4.16 7.1 ;
      RECT  0.98 7.1 4.16 96.64 ;
      RECT  4.16 3.7 447.74 4.16 ;
      RECT  4.16 7.1 447.74 96.64 ;
      RECT  447.74 3.7 450.92 4.16 ;
      RECT  447.74 4.16 450.92 7.1 ;
      RECT  447.74 7.1 450.92 96.64 ;
      RECT  0.98 396.74 4.16 435.96 ;
      RECT  0.98 435.96 4.16 438.9 ;
      RECT  0.98 438.9 4.16 439.36 ;
      RECT  4.16 396.74 447.74 435.96 ;
      RECT  4.16 438.9 447.74 439.36 ;
      RECT  447.74 396.74 450.92 435.96 ;
      RECT  447.74 435.96 450.92 438.9 ;
      RECT  447.74 438.9 450.92 439.36 ;
   LAYER  met4 ;
      RECT  86.44 0.98 88.02 442.44 ;
      RECT  88.02 0.62 92.56 0.98 ;
      RECT  94.14 0.62 98.0 0.98 ;
      RECT  99.58 0.62 103.44 0.98 ;
      RECT  105.02 0.62 109.56 0.98 ;
      RECT  111.14 0.62 115.0 0.98 ;
      RECT  116.58 0.62 121.8 0.98 ;
      RECT  64.22 0.62 69.44 0.98 ;
      RECT  71.02 0.62 74.88 0.98 ;
      RECT  88.02 0.98 381.56 442.08 ;
      RECT  381.56 0.98 383.14 442.08 ;
      RECT  377.7 442.08 381.56 442.44 ;
      RECT  372.26 442.08 376.12 442.44 ;
      RECT  76.46 0.62 80.32 0.98 ;
      RECT  81.9 0.62 86.44 0.98 ;
      RECT  123.38 0.62 124.52 0.98 ;
      RECT  126.1 0.62 126.56 0.98 ;
      RECT  128.14 0.62 150.36 0.98 ;
      RECT  151.94 0.62 175.52 0.98 ;
      RECT  177.1 0.62 200.68 0.98 ;
      RECT  202.26 0.62 225.84 0.98 ;
      RECT  227.42 0.62 250.32 0.98 ;
      RECT  251.9 0.62 275.48 0.98 ;
      RECT  277.06 0.62 300.64 0.98 ;
      RECT  88.02 442.08 125.88 442.44 ;
      RECT  127.46 442.08 151.04 442.44 ;
      RECT  152.62 442.08 176.2 442.44 ;
      RECT  177.78 442.08 201.36 442.44 ;
      RECT  202.94 442.08 225.84 442.44 ;
      RECT  227.42 442.08 250.32 442.44 ;
      RECT  251.9 442.08 276.16 442.44 ;
      RECT  277.74 442.08 301.32 442.44 ;
      RECT  302.9 442.08 370.68 442.44 ;
      RECT  451.14 0.98 451.28 442.08 ;
      RECT  383.14 442.08 448.2 442.3 ;
      RECT  383.14 442.3 448.2 442.44 ;
      RECT  448.2 442.3 451.14 442.44 ;
      RECT  451.14 442.08 451.28 442.3 ;
      RECT  451.14 442.3 451.28 442.44 ;
      RECT  302.22 0.62 448.2 0.76 ;
      RECT  302.22 0.76 448.2 0.98 ;
      RECT  448.2 0.62 451.14 0.76 ;
      RECT  451.14 0.62 451.28 0.76 ;
      RECT  451.14 0.76 451.28 0.98 ;
      RECT  0.62 0.98 0.76 442.3 ;
      RECT  0.62 442.3 0.76 442.44 ;
      RECT  0.76 442.3 3.7 442.44 ;
      RECT  3.7 442.3 86.44 442.44 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 0.98 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 62.64 0.76 ;
      RECT  3.7 0.76 62.64 0.98 ;
      RECT  3.7 0.98 4.16 4.16 ;
      RECT  3.7 4.16 4.16 438.9 ;
      RECT  3.7 438.9 4.16 442.3 ;
      RECT  4.16 0.98 7.1 4.16 ;
      RECT  4.16 438.9 7.1 442.3 ;
      RECT  7.1 0.98 86.44 4.16 ;
      RECT  7.1 4.16 86.44 438.9 ;
      RECT  7.1 438.9 86.44 442.3 ;
      RECT  383.14 0.98 444.8 4.16 ;
      RECT  383.14 4.16 444.8 438.9 ;
      RECT  383.14 438.9 444.8 442.08 ;
      RECT  444.8 0.98 447.74 4.16 ;
      RECT  444.8 438.9 447.74 442.08 ;
      RECT  447.74 0.98 448.2 4.16 ;
      RECT  447.74 4.16 448.2 438.9 ;
      RECT  447.74 438.9 448.2 442.08 ;
   END
END    sky130_sram_1kbyte_1rw1r_8x1024_8
END    LIBRARY
