**************************************************
* OpenRAM generated memory.
* Words: 512
* Data bits: 32
* Banks: 1
* Column mux: 4:1
* Trimmed: False
* LVS: False
**************************************************
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_cell_opt1.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_cell_opt1 BL BR VGND VPWR VPB VNB WL
X0 Q_bar WL BR VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
X1 Q Q_bar VGND VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
*X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
*X4 Q_bar WL Q_bar VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
X5 VPWR Q Q_bar VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X6 Q Q_bar VPWR VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X7 VGND Q Q_bar VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_cell_opt1a.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_cell_opt1a BL BR VGND VPWR VPB VNB WL
X0 Q_bar WL BR VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
X1 Q Q_bar VGND VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
*X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
*X4 Q_bar WL Q_bar VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
X5 VPWR Q Q_bar VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X6 Q Q_bar VPWR VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X7 VGND Q Q_bar VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_wlstrap.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_wlstrap VPWR
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_wlstrap_p.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_wlstrap_p VGND
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_wlstrapa.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_wlstrapa VPWR
.ends

.SUBCKT sky130_bitcell_array bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 vdd gnd
*.PININFO bl_0_0:B br_0_0:B bl_0_1:B br_0_1:B bl_0_2:B br_0_2:B bl_0_3:B br_0_3:B bl_0_4:B br_0_4:B bl_0_5:B br_0_5:B bl_0_6:B br_0_6:B bl_0_7:B br_0_7:B bl_0_8:B br_0_8:B bl_0_9:B br_0_9:B bl_0_10:B br_0_10:B bl_0_11:B br_0_11:B bl_0_12:B br_0_12:B bl_0_13:B br_0_13:B bl_0_14:B br_0_14:B bl_0_15:B br_0_15:B bl_0_16:B br_0_16:B bl_0_17:B br_0_17:B bl_0_18:B br_0_18:B bl_0_19:B br_0_19:B bl_0_20:B br_0_20:B bl_0_21:B br_0_21:B bl_0_22:B br_0_22:B bl_0_23:B br_0_23:B bl_0_24:B br_0_24:B bl_0_25:B br_0_25:B bl_0_26:B br_0_26:B bl_0_27:B br_0_27:B bl_0_28:B br_0_28:B bl_0_29:B br_0_29:B bl_0_30:B br_0_30:B bl_0_31:B br_0_31:B bl_0_32:B br_0_32:B bl_0_33:B br_0_33:B bl_0_34:B br_0_34:B bl_0_35:B br_0_35:B bl_0_36:B br_0_36:B bl_0_37:B br_0_37:B bl_0_38:B br_0_38:B bl_0_39:B br_0_39:B bl_0_40:B br_0_40:B bl_0_41:B br_0_41:B bl_0_42:B br_0_42:B bl_0_43:B br_0_43:B bl_0_44:B br_0_44:B bl_0_45:B br_0_45:B bl_0_46:B br_0_46:B bl_0_47:B br_0_47:B bl_0_48:B br_0_48:B bl_0_49:B br_0_49:B bl_0_50:B br_0_50:B bl_0_51:B br_0_51:B bl_0_52:B br_0_52:B bl_0_53:B br_0_53:B bl_0_54:B br_0_54:B bl_0_55:B br_0_55:B bl_0_56:B br_0_56:B bl_0_57:B br_0_57:B bl_0_58:B br_0_58:B bl_0_59:B br_0_59:B bl_0_60:B br_0_60:B bl_0_61:B br_0_61:B bl_0_62:B br_0_62:B bl_0_63:B br_0_63:B bl_0_64:B br_0_64:B bl_0_65:B br_0_65:B bl_0_66:B br_0_66:B bl_0_67:B br_0_67:B bl_0_68:B br_0_68:B bl_0_69:B br_0_69:B bl_0_70:B br_0_70:B bl_0_71:B br_0_71:B bl_0_72:B br_0_72:B bl_0_73:B br_0_73:B bl_0_74:B br_0_74:B bl_0_75:B br_0_75:B bl_0_76:B br_0_76:B bl_0_77:B br_0_77:B bl_0_78:B br_0_78:B bl_0_79:B br_0_79:B bl_0_80:B br_0_80:B bl_0_81:B br_0_81:B bl_0_82:B br_0_82:B bl_0_83:B br_0_83:B bl_0_84:B br_0_84:B bl_0_85:B br_0_85:B bl_0_86:B br_0_86:B bl_0_87:B br_0_87:B bl_0_88:B br_0_88:B bl_0_89:B br_0_89:B bl_0_90:B br_0_90:B bl_0_91:B br_0_91:B bl_0_92:B br_0_92:B bl_0_93:B br_0_93:B bl_0_94:B br_0_94:B bl_0_95:B br_0_95:B bl_0_96:B br_0_96:B bl_0_97:B br_0_97:B bl_0_98:B br_0_98:B bl_0_99:B br_0_99:B bl_0_100:B br_0_100:B bl_0_101:B br_0_101:B bl_0_102:B br_0_102:B bl_0_103:B br_0_103:B bl_0_104:B br_0_104:B bl_0_105:B br_0_105:B bl_0_106:B br_0_106:B bl_0_107:B br_0_107:B bl_0_108:B br_0_108:B bl_0_109:B br_0_109:B bl_0_110:B br_0_110:B bl_0_111:B br_0_111:B bl_0_112:B br_0_112:B bl_0_113:B br_0_113:B bl_0_114:B br_0_114:B bl_0_115:B br_0_115:B bl_0_116:B br_0_116:B bl_0_117:B br_0_117:B bl_0_118:B br_0_118:B bl_0_119:B br_0_119:B bl_0_120:B br_0_120:B bl_0_121:B br_0_121:B bl_0_122:B br_0_122:B bl_0_123:B br_0_123:B bl_0_124:B br_0_124:B bl_0_125:B br_0_125:B bl_0_126:B br_0_126:B bl_0_127:B br_0_127:B bl_0_128:B br_0_128:B wl_0_0:I wl_0_1:I wl_0_2:I wl_0_3:I wl_0_4:I wl_0_5:I wl_0_6:I wl_0_7:I wl_0_8:I wl_0_9:I wl_0_10:I wl_0_11:I wl_0_12:I wl_0_13:I wl_0_14:I wl_0_15:I wl_0_16:I wl_0_17:I wl_0_18:I wl_0_19:I wl_0_20:I wl_0_21:I wl_0_22:I wl_0_23:I wl_0_24:I wl_0_25:I wl_0_26:I wl_0_27:I wl_0_28:I wl_0_29:I wl_0_30:I wl_0_31:I wl_0_32:I wl_0_33:I wl_0_34:I wl_0_35:I wl_0_36:I wl_0_37:I wl_0_38:I wl_0_39:I wl_0_40:I wl_0_41:I wl_0_42:I wl_0_43:I wl_0_44:I wl_0_45:I wl_0_46:I wl_0_47:I wl_0_48:I wl_0_49:I wl_0_50:I wl_0_51:I wl_0_52:I wl_0_53:I wl_0_54:I wl_0_55:I wl_0_56:I wl_0_57:I wl_0_58:I wl_0_59:I wl_0_60:I wl_0_61:I wl_0_62:I wl_0_63:I wl_0_64:I wl_0_65:I wl_0_66:I wl_0_67:I wl_0_68:I wl_0_69:I wl_0_70:I wl_0_71:I wl_0_72:I wl_0_73:I wl_0_74:I wl_0_75:I wl_0_76:I wl_0_77:I wl_0_78:I wl_0_79:I wl_0_80:I wl_0_81:I wl_0_82:I wl_0_83:I wl_0_84:I wl_0_85:I wl_0_86:I wl_0_87:I wl_0_88:I wl_0_89:I wl_0_90:I wl_0_91:I wl_0_92:I wl_0_93:I wl_0_94:I wl_0_95:I wl_0_96:I wl_0_97:I wl_0_98:I wl_0_99:I wl_0_100:I wl_0_101:I wl_0_102:I wl_0_103:I wl_0_104:I wl_0_105:I wl_0_106:I wl_0_107:I wl_0_108:I wl_0_109:I wl_0_110:I wl_0_111:I wl_0_112:I wl_0_113:I wl_0_114:I wl_0_115:I wl_0_116:I wl_0_117:I wl_0_118:I wl_0_119:I wl_0_120:I wl_0_121:I wl_0_122:I wl_0_123:I wl_0_124:I wl_0_125:I wl_0_126:I wl_0_127:I wl_0_128:I vdd:B gnd:B
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* INPUT : wl_0_67 
* INPUT : wl_0_68 
* INPUT : wl_0_69 
* INPUT : wl_0_70 
* INPUT : wl_0_71 
* INPUT : wl_0_72 
* INPUT : wl_0_73 
* INPUT : wl_0_74 
* INPUT : wl_0_75 
* INPUT : wl_0_76 
* INPUT : wl_0_77 
* INPUT : wl_0_78 
* INPUT : wl_0_79 
* INPUT : wl_0_80 
* INPUT : wl_0_81 
* INPUT : wl_0_82 
* INPUT : wl_0_83 
* INPUT : wl_0_84 
* INPUT : wl_0_85 
* INPUT : wl_0_86 
* INPUT : wl_0_87 
* INPUT : wl_0_88 
* INPUT : wl_0_89 
* INPUT : wl_0_90 
* INPUT : wl_0_91 
* INPUT : wl_0_92 
* INPUT : wl_0_93 
* INPUT : wl_0_94 
* INPUT : wl_0_95 
* INPUT : wl_0_96 
* INPUT : wl_0_97 
* INPUT : wl_0_98 
* INPUT : wl_0_99 
* INPUT : wl_0_100 
* INPUT : wl_0_101 
* INPUT : wl_0_102 
* INPUT : wl_0_103 
* INPUT : wl_0_104 
* INPUT : wl_0_105 
* INPUT : wl_0_106 
* INPUT : wl_0_107 
* INPUT : wl_0_108 
* INPUT : wl_0_109 
* INPUT : wl_0_110 
* INPUT : wl_0_111 
* INPUT : wl_0_112 
* INPUT : wl_0_113 
* INPUT : wl_0_114 
* INPUT : wl_0_115 
* INPUT : wl_0_116 
* INPUT : wl_0_117 
* INPUT : wl_0_118 
* INPUT : wl_0_119 
* INPUT : wl_0_120 
* INPUT : wl_0_121 
* INPUT : wl_0_122 
* INPUT : wl_0_123 
* INPUT : wl_0_124 
* INPUT : wl_0_125 
* INPUT : wl_0_126 
* INPUT : wl_0_127 
* INPUT : wl_0_128 
* POWER : vdd 
* GROUND: gnd 
* rows: 129 cols: 129
Xrow_0_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_1_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_1_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_2_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_3_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_3_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_4_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_5_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_5_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_6_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_7_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_7_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_8_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_9_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_9_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_10_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_11_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_11_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_12_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_13_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_13_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_14_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_15_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_15_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_16_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_17_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_17_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_18_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_19_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_19_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_20_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_21_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_21_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_22_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_23_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_23_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_24_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_25_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_25_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_26_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_27_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_27_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_28_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_29_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_29_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_30_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_31_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_31_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_32_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_33_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_33_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_34_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_35_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_35_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_36_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_37_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_37_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_38_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_39_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_39_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_40_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_41_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_41_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_42_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_43_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_43_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_44_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_45_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_45_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_46_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_47_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_47_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_48_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_49_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_49_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_50_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_51_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_51_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_52_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_53_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_53_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_54_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_55_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_55_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_56_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_57_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_57_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_58_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_59_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_59_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_60_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_61_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_61_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_62_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_63_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_63_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_64_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_65_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_65_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_65_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_65_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_66_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_66_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_66_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_66_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_67_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_67_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_67_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_67_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_68_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_68_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_68_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_68_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_69_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_69_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_69_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_69_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_70_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_70_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_70_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_70_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_71_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_71_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_71_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_71_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_72_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_72_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_72_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_72_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_73_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_73_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_73_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_73_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_74_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_74_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_74_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_74_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_75_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_75_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_75_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_75_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_76_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_76_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_76_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_76_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_77_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_77_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_77_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_77_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_78_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_78_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_78_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_78_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_79_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_79_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_79_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_79_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_80_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_80_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_80_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_80_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_81_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_81_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_81_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_81_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_82_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_82_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_82_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_82_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_83_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_83_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_83_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_83_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_84_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_84_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_84_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_84_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_85_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_85_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_85_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_85_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_86_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_86_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_86_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_86_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_87_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_87_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_87_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_87_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_88_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_88_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_88_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_88_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_89_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_89_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_89_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_89_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_90_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_90_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_90_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_90_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_91_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_91_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_91_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_91_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_92_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_92_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_92_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_92_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_93_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_93_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_93_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_93_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_94_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_94_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_94_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_94_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_95_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_95_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_95_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_95_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_96_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_96_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_96_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_96_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_97_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_97_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_97_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_97_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_98_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_98_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_98_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_98_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_99_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_99_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_99_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_99_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_100_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_100_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_100_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_100_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_101_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_101_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_101_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_101_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_102_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_102_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_102_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_102_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_103_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_103_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_103_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_103_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_104_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_104_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_104_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_104_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_105_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_105_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_105_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_105_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_106_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_106_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_106_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_106_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_107_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_107_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_107_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_107_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_108_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_108_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_108_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_108_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_109_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_109_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_109_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_109_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_110_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_110_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_110_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_110_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_111_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_111_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_111_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_111_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_112_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_112_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_112_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_112_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_113_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_113_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_113_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_113_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_114_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_114_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_114_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_114_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_115_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_115_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_115_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_115_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_116_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_116_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_116_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_116_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_117_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_117_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_117_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_117_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_118_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_118_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_118_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_118_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_119_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_119_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_119_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_119_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_120_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_120_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_120_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_120_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_121_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_121_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_121_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_121_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_122_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_122_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_122_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_122_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_123_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_123_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_123_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_123_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_124_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_124_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_124_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_124_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_125_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_125_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_125_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_125_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_126_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_126_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_126_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_126_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_127_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_127_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_127_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_127_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_128_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_128_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_128_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_128_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__sram_sp_cell_opt1
.ENDS sky130_bitcell_array
* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_opt1_replica.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_cell_opt1_replica BL BR VGND VPWR VPB VNB WL
X0 VPWR WL BR VNB sky130_fd_pr__special_nfet_pass ad=4.375e+10p pd=920000u as=1.68e+10p ps=520000u w=140000u l=150000u
X1 Q VPWR VGND VNB sky130_fd_pr__special_nfet_latch ad=1.56e+11p pd=2.38e+06u as=8.08e+10p ps=1.28e+06u w=210000u l=150000u
X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass ad=1.68e+10p pd=520000u as=4.25e+10p ps=920000u w=140000u l=150000u
*X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass ad=3.5e+10p pd=780000u as=0p ps=0u w=70000u l=95000u
*X4 VPWR WL VPWR VPB sky130_fd_pr__special_pfet_pass ad=9.72e+10p pd=1.86e+06u as=0p ps=0u w=70000u l=95000u
X5 VPWR Q VPWR VPB sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X6 Q VPWR VPWR VPB sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X7 VGND Q VPWR VNB sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
.ends
* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_opt1a_replica.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_cell_opt1a_replica BL BR VGND VPWR VPB VNB WL
X0 VPWR WL BR VNB sky130_fd_pr__special_nfet_pass ad=4.375e+10p pd=920000u as=1.68e+10p ps=520000u w=140000u l=150000u
X1 Q VPWR VGND VNB sky130_fd_pr__special_nfet_latch ad=1.56e+11p pd=2.38e+06u as=8.08e+10p ps=1.28e+06u w=210000u l=150000u
X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass ad=1.68e+10p pd=520000u as=4.25e+10p ps=920000u w=140000u l=150000u
*X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass ad=3.5e+10p pd=780000u as=0p ps=0u w=70000u l=95000u
*X4 VPWR WL VPWR VPB sky130_fd_pr__special_pfet_pass ad=9.72e+10p pd=1.86e+06u as=0p ps=0u w=70000u l=95000u
X5 VPWR Q VPWR VPB sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X6 Q VPWR VPWR VPB sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X7 VGND Q VPWR VNB sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colend.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colend BL1 VPWR VGND BL0
*X0 BL1 a_0_24# BL1 w_96_0# sky130_fd_pr__nfet_01v8 ad=1.68e+10p pd=520000u as=0p ps=0u w=70000u l=210000u
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colenda.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colenda BL1 VPWR VGND BL0
*X0 BL1 a_0_24# BL1 w_96_0# sky130_fd_pr__nfet_01v8 ad=1.68e+10p pd=520000u as=0p ps=0u w=70000u l=210000u
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colend_p_cent.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colend_p_cent VGND VPB VNB
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colenda_p_cent.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colenda_p_cent VGND VPB VNB
.ends

.SUBCKT sky130_replica_column bl_0_0 br_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 wl_0_129 wl_0_130 wl_0_131 vdd gnd
*.PININFO bl_0_0:O br_0_0:O wl_0_0:I wl_0_1:I wl_0_2:I wl_0_3:I wl_0_4:I wl_0_5:I wl_0_6:I wl_0_7:I wl_0_8:I wl_0_9:I wl_0_10:I wl_0_11:I wl_0_12:I wl_0_13:I wl_0_14:I wl_0_15:I wl_0_16:I wl_0_17:I wl_0_18:I wl_0_19:I wl_0_20:I wl_0_21:I wl_0_22:I wl_0_23:I wl_0_24:I wl_0_25:I wl_0_26:I wl_0_27:I wl_0_28:I wl_0_29:I wl_0_30:I wl_0_31:I wl_0_32:I wl_0_33:I wl_0_34:I wl_0_35:I wl_0_36:I wl_0_37:I wl_0_38:I wl_0_39:I wl_0_40:I wl_0_41:I wl_0_42:I wl_0_43:I wl_0_44:I wl_0_45:I wl_0_46:I wl_0_47:I wl_0_48:I wl_0_49:I wl_0_50:I wl_0_51:I wl_0_52:I wl_0_53:I wl_0_54:I wl_0_55:I wl_0_56:I wl_0_57:I wl_0_58:I wl_0_59:I wl_0_60:I wl_0_61:I wl_0_62:I wl_0_63:I wl_0_64:I wl_0_65:I wl_0_66:I wl_0_67:I wl_0_68:I wl_0_69:I wl_0_70:I wl_0_71:I wl_0_72:I wl_0_73:I wl_0_74:I wl_0_75:I wl_0_76:I wl_0_77:I wl_0_78:I wl_0_79:I wl_0_80:I wl_0_81:I wl_0_82:I wl_0_83:I wl_0_84:I wl_0_85:I wl_0_86:I wl_0_87:I wl_0_88:I wl_0_89:I wl_0_90:I wl_0_91:I wl_0_92:I wl_0_93:I wl_0_94:I wl_0_95:I wl_0_96:I wl_0_97:I wl_0_98:I wl_0_99:I wl_0_100:I wl_0_101:I wl_0_102:I wl_0_103:I wl_0_104:I wl_0_105:I wl_0_106:I wl_0_107:I wl_0_108:I wl_0_109:I wl_0_110:I wl_0_111:I wl_0_112:I wl_0_113:I wl_0_114:I wl_0_115:I wl_0_116:I wl_0_117:I wl_0_118:I wl_0_119:I wl_0_120:I wl_0_121:I wl_0_122:I wl_0_123:I wl_0_124:I wl_0_125:I wl_0_126:I wl_0_127:I wl_0_128:I wl_0_129:I wl_0_130:I wl_0_131:I vdd:B gnd:B
* OUTPUT: bl_0_0 
* OUTPUT: br_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* INPUT : wl_0_67 
* INPUT : wl_0_68 
* INPUT : wl_0_69 
* INPUT : wl_0_70 
* INPUT : wl_0_71 
* INPUT : wl_0_72 
* INPUT : wl_0_73 
* INPUT : wl_0_74 
* INPUT : wl_0_75 
* INPUT : wl_0_76 
* INPUT : wl_0_77 
* INPUT : wl_0_78 
* INPUT : wl_0_79 
* INPUT : wl_0_80 
* INPUT : wl_0_81 
* INPUT : wl_0_82 
* INPUT : wl_0_83 
* INPUT : wl_0_84 
* INPUT : wl_0_85 
* INPUT : wl_0_86 
* INPUT : wl_0_87 
* INPUT : wl_0_88 
* INPUT : wl_0_89 
* INPUT : wl_0_90 
* INPUT : wl_0_91 
* INPUT : wl_0_92 
* INPUT : wl_0_93 
* INPUT : wl_0_94 
* INPUT : wl_0_95 
* INPUT : wl_0_96 
* INPUT : wl_0_97 
* INPUT : wl_0_98 
* INPUT : wl_0_99 
* INPUT : wl_0_100 
* INPUT : wl_0_101 
* INPUT : wl_0_102 
* INPUT : wl_0_103 
* INPUT : wl_0_104 
* INPUT : wl_0_105 
* INPUT : wl_0_106 
* INPUT : wl_0_107 
* INPUT : wl_0_108 
* INPUT : wl_0_109 
* INPUT : wl_0_110 
* INPUT : wl_0_111 
* INPUT : wl_0_112 
* INPUT : wl_0_113 
* INPUT : wl_0_114 
* INPUT : wl_0_115 
* INPUT : wl_0_116 
* INPUT : wl_0_117 
* INPUT : wl_0_118 
* INPUT : wl_0_119 
* INPUT : wl_0_120 
* INPUT : wl_0_121 
* INPUT : wl_0_122 
* INPUT : wl_0_123 
* INPUT : wl_0_124 
* INPUT : wl_0_125 
* INPUT : wl_0_126 
* INPUT : wl_0_127 
* INPUT : wl_0_128 
* INPUT : wl_0_129 
* INPUT : wl_0_130 
* INPUT : wl_0_131 
* POWER : vdd 
* GROUND: gnd 
Xrbc_0 bl_0_0 vdd gnd br_0_0 sky130_fd_bd_sram__sram_sp_colend
Xrbc_0_cap gnd gnd vdd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrbc_1 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_1 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_1_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_2 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_2 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_2_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_3 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_3 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_3_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_4 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_4 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_4_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_5 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_5 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_5_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_6 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_6 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_6_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_7 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_7 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_7_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_8 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_8 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_8_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_9 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_9 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_9_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_10 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_10 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_10_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_11 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_11 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_11_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_12 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_12 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_12_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_13 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_13 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_13_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_14 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_14 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_14_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_15 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_15 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_15_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_16 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_16 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_16_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_17 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_17 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_17_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_18 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_18 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_18_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_19 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_19 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_19_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_20 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_20 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_20_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_21 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_21 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_21_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_22 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_22 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_22_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_23 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_23 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_23_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_24 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_24 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_24_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_25 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_25 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_25_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_26 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_26 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_26_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_27 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_27 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_27_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_28 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_28 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_28_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_29 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_29 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_29_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_30 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_30 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_30_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_31 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_31 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_31_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_32 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_32 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_32_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_33 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_33 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_33_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_34 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_34 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_34_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_35 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_35 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_35_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_36 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_36 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_36_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_37 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_37 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_37_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_38 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_38 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_38_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_39 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_39 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_39_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_40 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_40 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_40_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_41 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_41 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_41_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_42 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_42 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_42_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_43 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_43 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_43_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_44 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_44 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_44_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_45 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_45 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_45_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_46 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_46 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_46_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_47 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_47 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_47_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_48 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_48 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_48_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_49 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_49 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_49_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_50 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_50 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_50_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_51 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_51 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_51_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_52 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_52 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_52_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_53 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_53 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_53_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_54 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_54 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_54_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_55 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_55 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_55_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_56 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_56 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_56_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_57 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_57 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_57_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_58 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_58 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_58_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_59 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_59 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_59_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_60 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_60 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_60_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_61 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_61 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_61_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_62 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_62 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_62_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_63 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_63 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_63_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_64 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_64 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_64_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_65 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_65 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_65_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_66 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_66 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_66_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_67 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_67 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_67_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_68 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_68 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_68_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_69 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_69 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_69_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_70 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_70 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_70_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_71 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_71 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_71_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_72 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_72 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_72_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_73 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_73 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_73_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_74 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_74 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_74_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_75 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_75 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_75_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_76 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_76 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_76_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_77 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_77 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_77_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_78 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_78 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_78_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_79 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_79 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_79_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_80 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_80 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_80_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_81 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_81 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_81_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_82 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_82 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_82_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_83 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_83 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_83_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_84 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_84 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_84_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_85 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_85 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_85_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_86 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_86 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_86_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_87 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_87 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_87_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_88 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_88 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_88_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_89 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_89 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_89_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_90 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_90 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_90_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_91 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_91 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_91_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_92 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_92 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_92_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_93 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_93 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_93_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_94 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_94 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_94_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_95 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_95 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_95_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_96 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_96 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_96_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_97 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_97 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_97_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_98 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_98 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_98_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_99 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_99 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_99_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_100 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_100 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_100_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_101 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_101 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_101_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_102 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_102 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_102_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_103 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_103 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_103_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_104 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_104 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_104_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_105 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_105 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_105_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_106 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_106 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_106_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_107 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_107 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_107_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_108 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_108 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_108_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_109 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_109 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_109_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_110 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_110 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_110_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_111 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_111 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_111_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_112 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_112 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_112_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_113 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_113 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_113_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_114 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_114 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_114_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_115 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_115 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_115_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_116 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_116 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_116_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_117 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_117 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_117_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_118 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_118 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_118_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_119 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_119 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_119_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_120 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_120 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_120_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_121 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_121 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_121_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_122 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_122 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_122_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_123 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_123 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_123_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_124 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_124 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_124_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_125 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_125 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_125_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_126 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_126 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_126_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_127 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_127 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_127_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_128 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_128 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_128_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_129 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_129 sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_129_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_130 bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_130 sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_130_strap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_131 bl_0_0 vdd gnd br_0_0 sky130_fd_bd_sram__sram_sp_colenda
Xrbc_131_cap gnd gnd vdd sky130_fd_bd_sram__sram_sp_colenda_p_cent
.ENDS sky130_replica_column
* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_opt1_dummy.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_cell_opt1_dummy BL BR VGND VPWR VPB VNB WL
X0 ll WL BR VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
X1 ul Q_bar_float VGND VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
X2 BL WL ul VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
*X3 ur WL ur VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
*X4 lr WL lr VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
X5 VPWR Q_float lr VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X6 ur Q_bar_float VPWR VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X7 VGND Q_float ll VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
.ends

* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy BL BR VGND VPWR VPB VNB WL
X0 ll WL BR VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
X1 ul Q_bar_float VGND VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
X2 BL WL ul VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
*X3 ur WL ur VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
*X4 lr WL lr VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
X5 VPWR Q_float lr VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X6 ur Q_bar_float VPWR VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X7 VGND Q_float ll VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
.ends

.SUBCKT sky130_dummy_array wl_0_0 dummy_bl_0 dummy_br_0 dummy_bl_1 dummy_br_1 dummy_bl_2 dummy_br_2 dummy_bl_3 dummy_br_3 dummy_bl_4 dummy_br_4 dummy_bl_5 dummy_br_5 dummy_bl_6 dummy_br_6 dummy_bl_7 dummy_br_7 dummy_bl_8 dummy_br_8 dummy_bl_9 dummy_br_9 dummy_bl_10 dummy_br_10 dummy_bl_11 dummy_br_11 dummy_bl_12 dummy_br_12 dummy_bl_13 dummy_br_13 dummy_bl_14 dummy_br_14 dummy_bl_15 dummy_br_15 dummy_bl_16 dummy_br_16 dummy_bl_17 dummy_br_17 dummy_bl_18 dummy_br_18 dummy_bl_19 dummy_br_19 dummy_bl_20 dummy_br_20 dummy_bl_21 dummy_br_21 dummy_bl_22 dummy_br_22 dummy_bl_23 dummy_br_23 dummy_bl_24 dummy_br_24 dummy_bl_25 dummy_br_25 dummy_bl_26 dummy_br_26 dummy_bl_27 dummy_br_27 dummy_bl_28 dummy_br_28 dummy_bl_29 dummy_br_29 dummy_bl_30 dummy_br_30 dummy_bl_31 dummy_br_31 dummy_bl_32 dummy_br_32 dummy_bl_33 dummy_br_33 dummy_bl_34 dummy_br_34 dummy_bl_35 dummy_br_35 dummy_bl_36 dummy_br_36 dummy_bl_37 dummy_br_37 dummy_bl_38 dummy_br_38 dummy_bl_39 dummy_br_39 dummy_bl_40 dummy_br_40 dummy_bl_41 dummy_br_41 dummy_bl_42 dummy_br_42 dummy_bl_43 dummy_br_43 dummy_bl_44 dummy_br_44 dummy_bl_45 dummy_br_45 dummy_bl_46 dummy_br_46 dummy_bl_47 dummy_br_47 dummy_bl_48 dummy_br_48 dummy_bl_49 dummy_br_49 dummy_bl_50 dummy_br_50 dummy_bl_51 dummy_br_51 dummy_bl_52 dummy_br_52 dummy_bl_53 dummy_br_53 dummy_bl_54 dummy_br_54 dummy_bl_55 dummy_br_55 dummy_bl_56 dummy_br_56 dummy_bl_57 dummy_br_57 dummy_bl_58 dummy_br_58 dummy_bl_59 dummy_br_59 dummy_bl_60 dummy_br_60 dummy_bl_61 dummy_br_61 dummy_bl_62 dummy_br_62 dummy_bl_63 dummy_br_63 dummy_bl_64 dummy_br_64 dummy_bl_65 dummy_br_65 dummy_bl_66 dummy_br_66 dummy_bl_67 dummy_br_67 dummy_bl_68 dummy_br_68 dummy_bl_69 dummy_br_69 dummy_bl_70 dummy_br_70 dummy_bl_71 dummy_br_71 dummy_bl_72 dummy_br_72 dummy_bl_73 dummy_br_73 dummy_bl_74 dummy_br_74 dummy_bl_75 dummy_br_75 dummy_bl_76 dummy_br_76 dummy_bl_77 dummy_br_77 dummy_bl_78 dummy_br_78 dummy_bl_79 dummy_br_79 dummy_bl_80 dummy_br_80 dummy_bl_81 dummy_br_81 dummy_bl_82 dummy_br_82 dummy_bl_83 dummy_br_83 dummy_bl_84 dummy_br_84 dummy_bl_85 dummy_br_85 dummy_bl_86 dummy_br_86 dummy_bl_87 dummy_br_87 dummy_bl_88 dummy_br_88 dummy_bl_89 dummy_br_89 dummy_bl_90 dummy_br_90 dummy_bl_91 dummy_br_91 dummy_bl_92 dummy_br_92 dummy_bl_93 dummy_br_93 dummy_bl_94 dummy_br_94 dummy_bl_95 dummy_br_95 dummy_bl_96 dummy_br_96 dummy_bl_97 dummy_br_97 dummy_bl_98 dummy_br_98 dummy_bl_99 dummy_br_99 dummy_bl_100 dummy_br_100 dummy_bl_101 dummy_br_101 dummy_bl_102 dummy_br_102 dummy_bl_103 dummy_br_103 dummy_bl_104 dummy_br_104 dummy_bl_105 dummy_br_105 dummy_bl_106 dummy_br_106 dummy_bl_107 dummy_br_107 dummy_bl_108 dummy_br_108 dummy_bl_109 dummy_br_109 dummy_bl_110 dummy_br_110 dummy_bl_111 dummy_br_111 dummy_bl_112 dummy_br_112 dummy_bl_113 dummy_br_113 dummy_bl_114 dummy_br_114 dummy_bl_115 dummy_br_115 dummy_bl_116 dummy_br_116 dummy_bl_117 dummy_br_117 dummy_bl_118 dummy_br_118 dummy_bl_119 dummy_br_119 dummy_bl_120 dummy_br_120 dummy_bl_121 dummy_br_121 dummy_bl_122 dummy_br_122 dummy_bl_123 dummy_br_123 dummy_bl_124 dummy_br_124 dummy_bl_125 dummy_br_125 dummy_bl_126 dummy_br_126 dummy_bl_127 dummy_br_127 dummy_bl_128 dummy_br_128 vdd gnd
*.PININFO wl_0_0:I dummy_bl_0:B dummy_br_0:B dummy_bl_1:B dummy_br_1:B dummy_bl_2:B dummy_br_2:B dummy_bl_3:B dummy_br_3:B dummy_bl_4:B dummy_br_4:B dummy_bl_5:B dummy_br_5:B dummy_bl_6:B dummy_br_6:B dummy_bl_7:B dummy_br_7:B dummy_bl_8:B dummy_br_8:B dummy_bl_9:B dummy_br_9:B dummy_bl_10:B dummy_br_10:B dummy_bl_11:B dummy_br_11:B dummy_bl_12:B dummy_br_12:B dummy_bl_13:B dummy_br_13:B dummy_bl_14:B dummy_br_14:B dummy_bl_15:B dummy_br_15:B dummy_bl_16:B dummy_br_16:B dummy_bl_17:B dummy_br_17:B dummy_bl_18:B dummy_br_18:B dummy_bl_19:B dummy_br_19:B dummy_bl_20:B dummy_br_20:B dummy_bl_21:B dummy_br_21:B dummy_bl_22:B dummy_br_22:B dummy_bl_23:B dummy_br_23:B dummy_bl_24:B dummy_br_24:B dummy_bl_25:B dummy_br_25:B dummy_bl_26:B dummy_br_26:B dummy_bl_27:B dummy_br_27:B dummy_bl_28:B dummy_br_28:B dummy_bl_29:B dummy_br_29:B dummy_bl_30:B dummy_br_30:B dummy_bl_31:B dummy_br_31:B dummy_bl_32:B dummy_br_32:B dummy_bl_33:B dummy_br_33:B dummy_bl_34:B dummy_br_34:B dummy_bl_35:B dummy_br_35:B dummy_bl_36:B dummy_br_36:B dummy_bl_37:B dummy_br_37:B dummy_bl_38:B dummy_br_38:B dummy_bl_39:B dummy_br_39:B dummy_bl_40:B dummy_br_40:B dummy_bl_41:B dummy_br_41:B dummy_bl_42:B dummy_br_42:B dummy_bl_43:B dummy_br_43:B dummy_bl_44:B dummy_br_44:B dummy_bl_45:B dummy_br_45:B dummy_bl_46:B dummy_br_46:B dummy_bl_47:B dummy_br_47:B dummy_bl_48:B dummy_br_48:B dummy_bl_49:B dummy_br_49:B dummy_bl_50:B dummy_br_50:B dummy_bl_51:B dummy_br_51:B dummy_bl_52:B dummy_br_52:B dummy_bl_53:B dummy_br_53:B dummy_bl_54:B dummy_br_54:B dummy_bl_55:B dummy_br_55:B dummy_bl_56:B dummy_br_56:B dummy_bl_57:B dummy_br_57:B dummy_bl_58:B dummy_br_58:B dummy_bl_59:B dummy_br_59:B dummy_bl_60:B dummy_br_60:B dummy_bl_61:B dummy_br_61:B dummy_bl_62:B dummy_br_62:B dummy_bl_63:B dummy_br_63:B dummy_bl_64:B dummy_br_64:B dummy_bl_65:B dummy_br_65:B dummy_bl_66:B dummy_br_66:B dummy_bl_67:B dummy_br_67:B dummy_bl_68:B dummy_br_68:B dummy_bl_69:B dummy_br_69:B dummy_bl_70:B dummy_br_70:B dummy_bl_71:B dummy_br_71:B dummy_bl_72:B dummy_br_72:B dummy_bl_73:B dummy_br_73:B dummy_bl_74:B dummy_br_74:B dummy_bl_75:B dummy_br_75:B dummy_bl_76:B dummy_br_76:B dummy_bl_77:B dummy_br_77:B dummy_bl_78:B dummy_br_78:B dummy_bl_79:B dummy_br_79:B dummy_bl_80:B dummy_br_80:B dummy_bl_81:B dummy_br_81:B dummy_bl_82:B dummy_br_82:B dummy_bl_83:B dummy_br_83:B dummy_bl_84:B dummy_br_84:B dummy_bl_85:B dummy_br_85:B dummy_bl_86:B dummy_br_86:B dummy_bl_87:B dummy_br_87:B dummy_bl_88:B dummy_br_88:B dummy_bl_89:B dummy_br_89:B dummy_bl_90:B dummy_br_90:B dummy_bl_91:B dummy_br_91:B dummy_bl_92:B dummy_br_92:B dummy_bl_93:B dummy_br_93:B dummy_bl_94:B dummy_br_94:B dummy_bl_95:B dummy_br_95:B dummy_bl_96:B dummy_br_96:B dummy_bl_97:B dummy_br_97:B dummy_bl_98:B dummy_br_98:B dummy_bl_99:B dummy_br_99:B dummy_bl_100:B dummy_br_100:B dummy_bl_101:B dummy_br_101:B dummy_bl_102:B dummy_br_102:B dummy_bl_103:B dummy_br_103:B dummy_bl_104:B dummy_br_104:B dummy_bl_105:B dummy_br_105:B dummy_bl_106:B dummy_br_106:B dummy_bl_107:B dummy_br_107:B dummy_bl_108:B dummy_br_108:B dummy_bl_109:B dummy_br_109:B dummy_bl_110:B dummy_br_110:B dummy_bl_111:B dummy_br_111:B dummy_bl_112:B dummy_br_112:B dummy_bl_113:B dummy_br_113:B dummy_bl_114:B dummy_br_114:B dummy_bl_115:B dummy_br_115:B dummy_bl_116:B dummy_br_116:B dummy_bl_117:B dummy_br_117:B dummy_bl_118:B dummy_br_118:B dummy_bl_119:B dummy_br_119:B dummy_bl_120:B dummy_br_120:B dummy_bl_121:B dummy_br_121:B dummy_bl_122:B dummy_br_122:B dummy_bl_123:B dummy_br_123:B dummy_bl_124:B dummy_br_124:B dummy_bl_125:B dummy_br_125:B dummy_bl_126:B dummy_br_126:B dummy_bl_127:B dummy_br_127:B dummy_bl_128:B dummy_br_128:B vdd:B gnd:B
* INPUT : wl_0_0 
* INOUT : dummy_bl_0 
* INOUT : dummy_br_0 
* INOUT : dummy_bl_1 
* INOUT : dummy_br_1 
* INOUT : dummy_bl_2 
* INOUT : dummy_br_2 
* INOUT : dummy_bl_3 
* INOUT : dummy_br_3 
* INOUT : dummy_bl_4 
* INOUT : dummy_br_4 
* INOUT : dummy_bl_5 
* INOUT : dummy_br_5 
* INOUT : dummy_bl_6 
* INOUT : dummy_br_6 
* INOUT : dummy_bl_7 
* INOUT : dummy_br_7 
* INOUT : dummy_bl_8 
* INOUT : dummy_br_8 
* INOUT : dummy_bl_9 
* INOUT : dummy_br_9 
* INOUT : dummy_bl_10 
* INOUT : dummy_br_10 
* INOUT : dummy_bl_11 
* INOUT : dummy_br_11 
* INOUT : dummy_bl_12 
* INOUT : dummy_br_12 
* INOUT : dummy_bl_13 
* INOUT : dummy_br_13 
* INOUT : dummy_bl_14 
* INOUT : dummy_br_14 
* INOUT : dummy_bl_15 
* INOUT : dummy_br_15 
* INOUT : dummy_bl_16 
* INOUT : dummy_br_16 
* INOUT : dummy_bl_17 
* INOUT : dummy_br_17 
* INOUT : dummy_bl_18 
* INOUT : dummy_br_18 
* INOUT : dummy_bl_19 
* INOUT : dummy_br_19 
* INOUT : dummy_bl_20 
* INOUT : dummy_br_20 
* INOUT : dummy_bl_21 
* INOUT : dummy_br_21 
* INOUT : dummy_bl_22 
* INOUT : dummy_br_22 
* INOUT : dummy_bl_23 
* INOUT : dummy_br_23 
* INOUT : dummy_bl_24 
* INOUT : dummy_br_24 
* INOUT : dummy_bl_25 
* INOUT : dummy_br_25 
* INOUT : dummy_bl_26 
* INOUT : dummy_br_26 
* INOUT : dummy_bl_27 
* INOUT : dummy_br_27 
* INOUT : dummy_bl_28 
* INOUT : dummy_br_28 
* INOUT : dummy_bl_29 
* INOUT : dummy_br_29 
* INOUT : dummy_bl_30 
* INOUT : dummy_br_30 
* INOUT : dummy_bl_31 
* INOUT : dummy_br_31 
* INOUT : dummy_bl_32 
* INOUT : dummy_br_32 
* INOUT : dummy_bl_33 
* INOUT : dummy_br_33 
* INOUT : dummy_bl_34 
* INOUT : dummy_br_34 
* INOUT : dummy_bl_35 
* INOUT : dummy_br_35 
* INOUT : dummy_bl_36 
* INOUT : dummy_br_36 
* INOUT : dummy_bl_37 
* INOUT : dummy_br_37 
* INOUT : dummy_bl_38 
* INOUT : dummy_br_38 
* INOUT : dummy_bl_39 
* INOUT : dummy_br_39 
* INOUT : dummy_bl_40 
* INOUT : dummy_br_40 
* INOUT : dummy_bl_41 
* INOUT : dummy_br_41 
* INOUT : dummy_bl_42 
* INOUT : dummy_br_42 
* INOUT : dummy_bl_43 
* INOUT : dummy_br_43 
* INOUT : dummy_bl_44 
* INOUT : dummy_br_44 
* INOUT : dummy_bl_45 
* INOUT : dummy_br_45 
* INOUT : dummy_bl_46 
* INOUT : dummy_br_46 
* INOUT : dummy_bl_47 
* INOUT : dummy_br_47 
* INOUT : dummy_bl_48 
* INOUT : dummy_br_48 
* INOUT : dummy_bl_49 
* INOUT : dummy_br_49 
* INOUT : dummy_bl_50 
* INOUT : dummy_br_50 
* INOUT : dummy_bl_51 
* INOUT : dummy_br_51 
* INOUT : dummy_bl_52 
* INOUT : dummy_br_52 
* INOUT : dummy_bl_53 
* INOUT : dummy_br_53 
* INOUT : dummy_bl_54 
* INOUT : dummy_br_54 
* INOUT : dummy_bl_55 
* INOUT : dummy_br_55 
* INOUT : dummy_bl_56 
* INOUT : dummy_br_56 
* INOUT : dummy_bl_57 
* INOUT : dummy_br_57 
* INOUT : dummy_bl_58 
* INOUT : dummy_br_58 
* INOUT : dummy_bl_59 
* INOUT : dummy_br_59 
* INOUT : dummy_bl_60 
* INOUT : dummy_br_60 
* INOUT : dummy_bl_61 
* INOUT : dummy_br_61 
* INOUT : dummy_bl_62 
* INOUT : dummy_br_62 
* INOUT : dummy_bl_63 
* INOUT : dummy_br_63 
* INOUT : dummy_bl_64 
* INOUT : dummy_br_64 
* INOUT : dummy_bl_65 
* INOUT : dummy_br_65 
* INOUT : dummy_bl_66 
* INOUT : dummy_br_66 
* INOUT : dummy_bl_67 
* INOUT : dummy_br_67 
* INOUT : dummy_bl_68 
* INOUT : dummy_br_68 
* INOUT : dummy_bl_69 
* INOUT : dummy_br_69 
* INOUT : dummy_bl_70 
* INOUT : dummy_br_70 
* INOUT : dummy_bl_71 
* INOUT : dummy_br_71 
* INOUT : dummy_bl_72 
* INOUT : dummy_br_72 
* INOUT : dummy_bl_73 
* INOUT : dummy_br_73 
* INOUT : dummy_bl_74 
* INOUT : dummy_br_74 
* INOUT : dummy_bl_75 
* INOUT : dummy_br_75 
* INOUT : dummy_bl_76 
* INOUT : dummy_br_76 
* INOUT : dummy_bl_77 
* INOUT : dummy_br_77 
* INOUT : dummy_bl_78 
* INOUT : dummy_br_78 
* INOUT : dummy_bl_79 
* INOUT : dummy_br_79 
* INOUT : dummy_bl_80 
* INOUT : dummy_br_80 
* INOUT : dummy_bl_81 
* INOUT : dummy_br_81 
* INOUT : dummy_bl_82 
* INOUT : dummy_br_82 
* INOUT : dummy_bl_83 
* INOUT : dummy_br_83 
* INOUT : dummy_bl_84 
* INOUT : dummy_br_84 
* INOUT : dummy_bl_85 
* INOUT : dummy_br_85 
* INOUT : dummy_bl_86 
* INOUT : dummy_br_86 
* INOUT : dummy_bl_87 
* INOUT : dummy_br_87 
* INOUT : dummy_bl_88 
* INOUT : dummy_br_88 
* INOUT : dummy_bl_89 
* INOUT : dummy_br_89 
* INOUT : dummy_bl_90 
* INOUT : dummy_br_90 
* INOUT : dummy_bl_91 
* INOUT : dummy_br_91 
* INOUT : dummy_bl_92 
* INOUT : dummy_br_92 
* INOUT : dummy_bl_93 
* INOUT : dummy_br_93 
* INOUT : dummy_bl_94 
* INOUT : dummy_br_94 
* INOUT : dummy_bl_95 
* INOUT : dummy_br_95 
* INOUT : dummy_bl_96 
* INOUT : dummy_br_96 
* INOUT : dummy_bl_97 
* INOUT : dummy_br_97 
* INOUT : dummy_bl_98 
* INOUT : dummy_br_98 
* INOUT : dummy_bl_99 
* INOUT : dummy_br_99 
* INOUT : dummy_bl_100 
* INOUT : dummy_br_100 
* INOUT : dummy_bl_101 
* INOUT : dummy_br_101 
* INOUT : dummy_bl_102 
* INOUT : dummy_br_102 
* INOUT : dummy_bl_103 
* INOUT : dummy_br_103 
* INOUT : dummy_bl_104 
* INOUT : dummy_br_104 
* INOUT : dummy_bl_105 
* INOUT : dummy_br_105 
* INOUT : dummy_bl_106 
* INOUT : dummy_br_106 
* INOUT : dummy_bl_107 
* INOUT : dummy_br_107 
* INOUT : dummy_bl_108 
* INOUT : dummy_br_108 
* INOUT : dummy_bl_109 
* INOUT : dummy_br_109 
* INOUT : dummy_bl_110 
* INOUT : dummy_br_110 
* INOUT : dummy_bl_111 
* INOUT : dummy_br_111 
* INOUT : dummy_bl_112 
* INOUT : dummy_br_112 
* INOUT : dummy_bl_113 
* INOUT : dummy_br_113 
* INOUT : dummy_bl_114 
* INOUT : dummy_br_114 
* INOUT : dummy_bl_115 
* INOUT : dummy_br_115 
* INOUT : dummy_bl_116 
* INOUT : dummy_br_116 
* INOUT : dummy_bl_117 
* INOUT : dummy_br_117 
* INOUT : dummy_bl_118 
* INOUT : dummy_br_118 
* INOUT : dummy_bl_119 
* INOUT : dummy_br_119 
* INOUT : dummy_bl_120 
* INOUT : dummy_br_120 
* INOUT : dummy_bl_121 
* INOUT : dummy_br_121 
* INOUT : dummy_bl_122 
* INOUT : dummy_br_122 
* INOUT : dummy_bl_123 
* INOUT : dummy_br_123 
* INOUT : dummy_bl_124 
* INOUT : dummy_br_124 
* INOUT : dummy_bl_125 
* INOUT : dummy_br_125 
* INOUT : dummy_bl_126 
* INOUT : dummy_br_126 
* INOUT : dummy_bl_127 
* INOUT : dummy_br_127 
* INOUT : dummy_bl_128 
* INOUT : dummy_br_128 
* POWER : vdd 
* GROUND: gnd 
Xrow_0_col_0_bitcell bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_0_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_1_bitcell bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_1_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_2_bitcell bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_2_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_3_bitcell bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_3_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_4_bitcell bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_4_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_5_bitcell bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_5_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_6_bitcell bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_6_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_7_bitcell bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_7_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_8_bitcell bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_8_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_9_bitcell bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_9_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_10_bitcell bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_10_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_11_bitcell bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_11_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_12_bitcell bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_12_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_13_bitcell bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_13_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_14_bitcell bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_14_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_15_bitcell bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_15_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_16_bitcell bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_16_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_17_bitcell bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_17_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_18_bitcell bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_18_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_19_bitcell bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_19_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_20_bitcell bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_20_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_21_bitcell bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_21_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_22_bitcell bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_22_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_23_bitcell bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_23_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_24_bitcell bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_24_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_25_bitcell bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_25_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_26_bitcell bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_26_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_27_bitcell bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_27_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_28_bitcell bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_28_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_29_bitcell bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_29_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_30_bitcell bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_30_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_31_bitcell bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_31_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_32_bitcell bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_32_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_33_bitcell bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_33_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_34_bitcell bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_34_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_35_bitcell bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_35_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_36_bitcell bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_36_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_37_bitcell bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_37_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_38_bitcell bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_38_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_39_bitcell bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_39_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_40_bitcell bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_40_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_41_bitcell bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_41_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_42_bitcell bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_42_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_43_bitcell bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_43_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_44_bitcell bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_44_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_45_bitcell bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_45_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_46_bitcell bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_46_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_47_bitcell bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_47_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_48_bitcell bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_48_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_49_bitcell bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_49_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_50_bitcell bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_50_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_51_bitcell bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_51_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_52_bitcell bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_52_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_53_bitcell bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_53_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_54_bitcell bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_54_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_55_bitcell bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_55_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_56_bitcell bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_56_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_57_bitcell bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_57_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_58_bitcell bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_58_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_59_bitcell bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_59_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_60_bitcell bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_60_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_61_bitcell bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_61_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_62_bitcell bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_62_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_63_bitcell bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_63_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_64_bitcell bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_64_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_65_bitcell bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_65_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_66_bitcell bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_66_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_67_bitcell bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_67_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_68_bitcell bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_68_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_69_bitcell bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_69_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_70_bitcell bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_70_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_71_bitcell bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_71_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_72_bitcell bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_72_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_73_bitcell bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_73_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_74_bitcell bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_74_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_75_bitcell bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_75_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_76_bitcell bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_76_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_77_bitcell bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_77_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_78_bitcell bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_78_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_79_bitcell bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_79_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_80_bitcell bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_80_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_81_bitcell bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_81_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_82_bitcell bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_82_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_83_bitcell bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_83_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_84_bitcell bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_84_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_85_bitcell bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_85_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_86_bitcell bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_86_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_87_bitcell bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_87_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_88_bitcell bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_88_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_89_bitcell bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_89_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_90_bitcell bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_90_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_91_bitcell bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_91_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_92_bitcell bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_92_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_93_bitcell bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_93_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_94_bitcell bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_94_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_95_bitcell bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_95_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_96_bitcell bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_96_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_97_bitcell bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_97_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_98_bitcell bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_98_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_99_bitcell bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_99_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_100_bitcell bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_100_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_101_bitcell bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_101_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_102_bitcell bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_102_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_103_bitcell bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_103_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_104_bitcell bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_104_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_105_bitcell bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_105_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_106_bitcell bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_106_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_107_bitcell bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_107_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_108_bitcell bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_108_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_109_bitcell bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_109_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_110_bitcell bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_110_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_111_bitcell bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_111_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_112_bitcell bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_112_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_113_bitcell bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_113_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_114_bitcell bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_114_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_115_bitcell bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_115_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_116_bitcell bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_116_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_117_bitcell bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_117_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_118_bitcell bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_118_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_119_bitcell bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_119_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_120_bitcell bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_120_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_121_bitcell bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_121_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_122_bitcell bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_122_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_123_bitcell bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_123_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_124_bitcell bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_124_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_125_bitcell bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_125_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_126_bitcell bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_126_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_127_bitcell bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_127_wlstrap vdd sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_128_bitcell bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_0 sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
.ENDS sky130_dummy_array
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colend_cent.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colend_cent VPWR VPB VNB
.ends

.SUBCKT sky130_col_cap_array fake_bl_0 fake_br_0 fake_bl_1 fake_br_1 fake_bl_2 fake_br_2 fake_bl_3 fake_br_3 fake_bl_4 fake_br_4 fake_bl_5 fake_br_5 fake_bl_6 fake_br_6 fake_bl_7 fake_br_7 fake_bl_8 fake_br_8 fake_bl_9 fake_br_9 fake_bl_10 fake_br_10 fake_bl_11 fake_br_11 fake_bl_12 fake_br_12 fake_bl_13 fake_br_13 fake_bl_14 fake_br_14 fake_bl_15 fake_br_15 fake_bl_16 fake_br_16 fake_bl_17 fake_br_17 fake_bl_18 fake_br_18 fake_bl_19 fake_br_19 fake_bl_20 fake_br_20 fake_bl_21 fake_br_21 fake_bl_22 fake_br_22 fake_bl_23 fake_br_23 fake_bl_24 fake_br_24 fake_bl_25 fake_br_25 fake_bl_26 fake_br_26 fake_bl_27 fake_br_27 fake_bl_28 fake_br_28 fake_bl_29 fake_br_29 fake_bl_30 fake_br_30 fake_bl_31 fake_br_31 fake_bl_32 fake_br_32 fake_bl_33 fake_br_33 fake_bl_34 fake_br_34 fake_bl_35 fake_br_35 fake_bl_36 fake_br_36 fake_bl_37 fake_br_37 fake_bl_38 fake_br_38 fake_bl_39 fake_br_39 fake_bl_40 fake_br_40 fake_bl_41 fake_br_41 fake_bl_42 fake_br_42 fake_bl_43 fake_br_43 fake_bl_44 fake_br_44 fake_bl_45 fake_br_45 fake_bl_46 fake_br_46 fake_bl_47 fake_br_47 fake_bl_48 fake_br_48 fake_bl_49 fake_br_49 fake_bl_50 fake_br_50 fake_bl_51 fake_br_51 fake_bl_52 fake_br_52 fake_bl_53 fake_br_53 fake_bl_54 fake_br_54 fake_bl_55 fake_br_55 fake_bl_56 fake_br_56 fake_bl_57 fake_br_57 fake_bl_58 fake_br_58 fake_bl_59 fake_br_59 fake_bl_60 fake_br_60 fake_bl_61 fake_br_61 fake_bl_62 fake_br_62 fake_bl_63 fake_br_63 fake_bl_64 fake_br_64 fake_bl_65 fake_br_65 fake_bl_66 fake_br_66 fake_bl_67 fake_br_67 fake_bl_68 fake_br_68 fake_bl_69 fake_br_69 fake_bl_70 fake_br_70 fake_bl_71 fake_br_71 fake_bl_72 fake_br_72 fake_bl_73 fake_br_73 fake_bl_74 fake_br_74 fake_bl_75 fake_br_75 fake_bl_76 fake_br_76 fake_bl_77 fake_br_77 fake_bl_78 fake_br_78 fake_bl_79 fake_br_79 fake_bl_80 fake_br_80 fake_bl_81 fake_br_81 fake_bl_82 fake_br_82 fake_bl_83 fake_br_83 fake_bl_84 fake_br_84 fake_bl_85 fake_br_85 fake_bl_86 fake_br_86 fake_bl_87 fake_br_87 fake_bl_88 fake_br_88 fake_bl_89 fake_br_89 fake_bl_90 fake_br_90 fake_bl_91 fake_br_91 fake_bl_92 fake_br_92 fake_bl_93 fake_br_93 fake_bl_94 fake_br_94 fake_bl_95 fake_br_95 fake_bl_96 fake_br_96 fake_bl_97 fake_br_97 fake_bl_98 fake_br_98 fake_bl_99 fake_br_99 fake_bl_100 fake_br_100 fake_bl_101 fake_br_101 fake_bl_102 fake_br_102 fake_bl_103 fake_br_103 fake_bl_104 fake_br_104 fake_bl_105 fake_br_105 fake_bl_106 fake_br_106 fake_bl_107 fake_br_107 fake_bl_108 fake_br_108 fake_bl_109 fake_br_109 fake_bl_110 fake_br_110 fake_bl_111 fake_br_111 fake_bl_112 fake_br_112 fake_bl_113 fake_br_113 fake_bl_114 fake_br_114 fake_bl_115 fake_br_115 fake_bl_116 fake_br_116 fake_bl_117 fake_br_117 fake_bl_118 fake_br_118 fake_bl_119 fake_br_119 fake_bl_120 fake_br_120 fake_bl_121 fake_br_121 fake_bl_122 fake_br_122 fake_bl_123 fake_br_123 fake_bl_124 fake_br_124 fake_bl_125 fake_br_125 fake_bl_126 fake_br_126 fake_bl_127 fake_br_127 fake_bl_128 fake_br_128 fake_wl vdd gnd
*.PININFO fake_bl_0:O fake_br_0:O fake_bl_1:O fake_br_1:O fake_bl_2:O fake_br_2:O fake_bl_3:O fake_br_3:O fake_bl_4:O fake_br_4:O fake_bl_5:O fake_br_5:O fake_bl_6:O fake_br_6:O fake_bl_7:O fake_br_7:O fake_bl_8:O fake_br_8:O fake_bl_9:O fake_br_9:O fake_bl_10:O fake_br_10:O fake_bl_11:O fake_br_11:O fake_bl_12:O fake_br_12:O fake_bl_13:O fake_br_13:O fake_bl_14:O fake_br_14:O fake_bl_15:O fake_br_15:O fake_bl_16:O fake_br_16:O fake_bl_17:O fake_br_17:O fake_bl_18:O fake_br_18:O fake_bl_19:O fake_br_19:O fake_bl_20:O fake_br_20:O fake_bl_21:O fake_br_21:O fake_bl_22:O fake_br_22:O fake_bl_23:O fake_br_23:O fake_bl_24:O fake_br_24:O fake_bl_25:O fake_br_25:O fake_bl_26:O fake_br_26:O fake_bl_27:O fake_br_27:O fake_bl_28:O fake_br_28:O fake_bl_29:O fake_br_29:O fake_bl_30:O fake_br_30:O fake_bl_31:O fake_br_31:O fake_bl_32:O fake_br_32:O fake_bl_33:O fake_br_33:O fake_bl_34:O fake_br_34:O fake_bl_35:O fake_br_35:O fake_bl_36:O fake_br_36:O fake_bl_37:O fake_br_37:O fake_bl_38:O fake_br_38:O fake_bl_39:O fake_br_39:O fake_bl_40:O fake_br_40:O fake_bl_41:O fake_br_41:O fake_bl_42:O fake_br_42:O fake_bl_43:O fake_br_43:O fake_bl_44:O fake_br_44:O fake_bl_45:O fake_br_45:O fake_bl_46:O fake_br_46:O fake_bl_47:O fake_br_47:O fake_bl_48:O fake_br_48:O fake_bl_49:O fake_br_49:O fake_bl_50:O fake_br_50:O fake_bl_51:O fake_br_51:O fake_bl_52:O fake_br_52:O fake_bl_53:O fake_br_53:O fake_bl_54:O fake_br_54:O fake_bl_55:O fake_br_55:O fake_bl_56:O fake_br_56:O fake_bl_57:O fake_br_57:O fake_bl_58:O fake_br_58:O fake_bl_59:O fake_br_59:O fake_bl_60:O fake_br_60:O fake_bl_61:O fake_br_61:O fake_bl_62:O fake_br_62:O fake_bl_63:O fake_br_63:O fake_bl_64:O fake_br_64:O fake_bl_65:O fake_br_65:O fake_bl_66:O fake_br_66:O fake_bl_67:O fake_br_67:O fake_bl_68:O fake_br_68:O fake_bl_69:O fake_br_69:O fake_bl_70:O fake_br_70:O fake_bl_71:O fake_br_71:O fake_bl_72:O fake_br_72:O fake_bl_73:O fake_br_73:O fake_bl_74:O fake_br_74:O fake_bl_75:O fake_br_75:O fake_bl_76:O fake_br_76:O fake_bl_77:O fake_br_77:O fake_bl_78:O fake_br_78:O fake_bl_79:O fake_br_79:O fake_bl_80:O fake_br_80:O fake_bl_81:O fake_br_81:O fake_bl_82:O fake_br_82:O fake_bl_83:O fake_br_83:O fake_bl_84:O fake_br_84:O fake_bl_85:O fake_br_85:O fake_bl_86:O fake_br_86:O fake_bl_87:O fake_br_87:O fake_bl_88:O fake_br_88:O fake_bl_89:O fake_br_89:O fake_bl_90:O fake_br_90:O fake_bl_91:O fake_br_91:O fake_bl_92:O fake_br_92:O fake_bl_93:O fake_br_93:O fake_bl_94:O fake_br_94:O fake_bl_95:O fake_br_95:O fake_bl_96:O fake_br_96:O fake_bl_97:O fake_br_97:O fake_bl_98:O fake_br_98:O fake_bl_99:O fake_br_99:O fake_bl_100:O fake_br_100:O fake_bl_101:O fake_br_101:O fake_bl_102:O fake_br_102:O fake_bl_103:O fake_br_103:O fake_bl_104:O fake_br_104:O fake_bl_105:O fake_br_105:O fake_bl_106:O fake_br_106:O fake_bl_107:O fake_br_107:O fake_bl_108:O fake_br_108:O fake_bl_109:O fake_br_109:O fake_bl_110:O fake_br_110:O fake_bl_111:O fake_br_111:O fake_bl_112:O fake_br_112:O fake_bl_113:O fake_br_113:O fake_bl_114:O fake_br_114:O fake_bl_115:O fake_br_115:O fake_bl_116:O fake_br_116:O fake_bl_117:O fake_br_117:O fake_bl_118:O fake_br_118:O fake_bl_119:O fake_br_119:O fake_bl_120:O fake_br_120:O fake_bl_121:O fake_br_121:O fake_bl_122:O fake_br_122:O fake_bl_123:O fake_br_123:O fake_bl_124:O fake_br_124:O fake_bl_125:O fake_br_125:O fake_bl_126:O fake_br_126:O fake_bl_127:O fake_br_127:O fake_bl_128:O fake_br_128:O fake_wl:I vdd:B gnd:B
* OUTPUT: fake_bl_0 
* OUTPUT: fake_br_0 
* OUTPUT: fake_bl_1 
* OUTPUT: fake_br_1 
* OUTPUT: fake_bl_2 
* OUTPUT: fake_br_2 
* OUTPUT: fake_bl_3 
* OUTPUT: fake_br_3 
* OUTPUT: fake_bl_4 
* OUTPUT: fake_br_4 
* OUTPUT: fake_bl_5 
* OUTPUT: fake_br_5 
* OUTPUT: fake_bl_6 
* OUTPUT: fake_br_6 
* OUTPUT: fake_bl_7 
* OUTPUT: fake_br_7 
* OUTPUT: fake_bl_8 
* OUTPUT: fake_br_8 
* OUTPUT: fake_bl_9 
* OUTPUT: fake_br_9 
* OUTPUT: fake_bl_10 
* OUTPUT: fake_br_10 
* OUTPUT: fake_bl_11 
* OUTPUT: fake_br_11 
* OUTPUT: fake_bl_12 
* OUTPUT: fake_br_12 
* OUTPUT: fake_bl_13 
* OUTPUT: fake_br_13 
* OUTPUT: fake_bl_14 
* OUTPUT: fake_br_14 
* OUTPUT: fake_bl_15 
* OUTPUT: fake_br_15 
* OUTPUT: fake_bl_16 
* OUTPUT: fake_br_16 
* OUTPUT: fake_bl_17 
* OUTPUT: fake_br_17 
* OUTPUT: fake_bl_18 
* OUTPUT: fake_br_18 
* OUTPUT: fake_bl_19 
* OUTPUT: fake_br_19 
* OUTPUT: fake_bl_20 
* OUTPUT: fake_br_20 
* OUTPUT: fake_bl_21 
* OUTPUT: fake_br_21 
* OUTPUT: fake_bl_22 
* OUTPUT: fake_br_22 
* OUTPUT: fake_bl_23 
* OUTPUT: fake_br_23 
* OUTPUT: fake_bl_24 
* OUTPUT: fake_br_24 
* OUTPUT: fake_bl_25 
* OUTPUT: fake_br_25 
* OUTPUT: fake_bl_26 
* OUTPUT: fake_br_26 
* OUTPUT: fake_bl_27 
* OUTPUT: fake_br_27 
* OUTPUT: fake_bl_28 
* OUTPUT: fake_br_28 
* OUTPUT: fake_bl_29 
* OUTPUT: fake_br_29 
* OUTPUT: fake_bl_30 
* OUTPUT: fake_br_30 
* OUTPUT: fake_bl_31 
* OUTPUT: fake_br_31 
* OUTPUT: fake_bl_32 
* OUTPUT: fake_br_32 
* OUTPUT: fake_bl_33 
* OUTPUT: fake_br_33 
* OUTPUT: fake_bl_34 
* OUTPUT: fake_br_34 
* OUTPUT: fake_bl_35 
* OUTPUT: fake_br_35 
* OUTPUT: fake_bl_36 
* OUTPUT: fake_br_36 
* OUTPUT: fake_bl_37 
* OUTPUT: fake_br_37 
* OUTPUT: fake_bl_38 
* OUTPUT: fake_br_38 
* OUTPUT: fake_bl_39 
* OUTPUT: fake_br_39 
* OUTPUT: fake_bl_40 
* OUTPUT: fake_br_40 
* OUTPUT: fake_bl_41 
* OUTPUT: fake_br_41 
* OUTPUT: fake_bl_42 
* OUTPUT: fake_br_42 
* OUTPUT: fake_bl_43 
* OUTPUT: fake_br_43 
* OUTPUT: fake_bl_44 
* OUTPUT: fake_br_44 
* OUTPUT: fake_bl_45 
* OUTPUT: fake_br_45 
* OUTPUT: fake_bl_46 
* OUTPUT: fake_br_46 
* OUTPUT: fake_bl_47 
* OUTPUT: fake_br_47 
* OUTPUT: fake_bl_48 
* OUTPUT: fake_br_48 
* OUTPUT: fake_bl_49 
* OUTPUT: fake_br_49 
* OUTPUT: fake_bl_50 
* OUTPUT: fake_br_50 
* OUTPUT: fake_bl_51 
* OUTPUT: fake_br_51 
* OUTPUT: fake_bl_52 
* OUTPUT: fake_br_52 
* OUTPUT: fake_bl_53 
* OUTPUT: fake_br_53 
* OUTPUT: fake_bl_54 
* OUTPUT: fake_br_54 
* OUTPUT: fake_bl_55 
* OUTPUT: fake_br_55 
* OUTPUT: fake_bl_56 
* OUTPUT: fake_br_56 
* OUTPUT: fake_bl_57 
* OUTPUT: fake_br_57 
* OUTPUT: fake_bl_58 
* OUTPUT: fake_br_58 
* OUTPUT: fake_bl_59 
* OUTPUT: fake_br_59 
* OUTPUT: fake_bl_60 
* OUTPUT: fake_br_60 
* OUTPUT: fake_bl_61 
* OUTPUT: fake_br_61 
* OUTPUT: fake_bl_62 
* OUTPUT: fake_br_62 
* OUTPUT: fake_bl_63 
* OUTPUT: fake_br_63 
* OUTPUT: fake_bl_64 
* OUTPUT: fake_br_64 
* OUTPUT: fake_bl_65 
* OUTPUT: fake_br_65 
* OUTPUT: fake_bl_66 
* OUTPUT: fake_br_66 
* OUTPUT: fake_bl_67 
* OUTPUT: fake_br_67 
* OUTPUT: fake_bl_68 
* OUTPUT: fake_br_68 
* OUTPUT: fake_bl_69 
* OUTPUT: fake_br_69 
* OUTPUT: fake_bl_70 
* OUTPUT: fake_br_70 
* OUTPUT: fake_bl_71 
* OUTPUT: fake_br_71 
* OUTPUT: fake_bl_72 
* OUTPUT: fake_br_72 
* OUTPUT: fake_bl_73 
* OUTPUT: fake_br_73 
* OUTPUT: fake_bl_74 
* OUTPUT: fake_br_74 
* OUTPUT: fake_bl_75 
* OUTPUT: fake_br_75 
* OUTPUT: fake_bl_76 
* OUTPUT: fake_br_76 
* OUTPUT: fake_bl_77 
* OUTPUT: fake_br_77 
* OUTPUT: fake_bl_78 
* OUTPUT: fake_br_78 
* OUTPUT: fake_bl_79 
* OUTPUT: fake_br_79 
* OUTPUT: fake_bl_80 
* OUTPUT: fake_br_80 
* OUTPUT: fake_bl_81 
* OUTPUT: fake_br_81 
* OUTPUT: fake_bl_82 
* OUTPUT: fake_br_82 
* OUTPUT: fake_bl_83 
* OUTPUT: fake_br_83 
* OUTPUT: fake_bl_84 
* OUTPUT: fake_br_84 
* OUTPUT: fake_bl_85 
* OUTPUT: fake_br_85 
* OUTPUT: fake_bl_86 
* OUTPUT: fake_br_86 
* OUTPUT: fake_bl_87 
* OUTPUT: fake_br_87 
* OUTPUT: fake_bl_88 
* OUTPUT: fake_br_88 
* OUTPUT: fake_bl_89 
* OUTPUT: fake_br_89 
* OUTPUT: fake_bl_90 
* OUTPUT: fake_br_90 
* OUTPUT: fake_bl_91 
* OUTPUT: fake_br_91 
* OUTPUT: fake_bl_92 
* OUTPUT: fake_br_92 
* OUTPUT: fake_bl_93 
* OUTPUT: fake_br_93 
* OUTPUT: fake_bl_94 
* OUTPUT: fake_br_94 
* OUTPUT: fake_bl_95 
* OUTPUT: fake_br_95 
* OUTPUT: fake_bl_96 
* OUTPUT: fake_br_96 
* OUTPUT: fake_bl_97 
* OUTPUT: fake_br_97 
* OUTPUT: fake_bl_98 
* OUTPUT: fake_br_98 
* OUTPUT: fake_bl_99 
* OUTPUT: fake_br_99 
* OUTPUT: fake_bl_100 
* OUTPUT: fake_br_100 
* OUTPUT: fake_bl_101 
* OUTPUT: fake_br_101 
* OUTPUT: fake_bl_102 
* OUTPUT: fake_br_102 
* OUTPUT: fake_bl_103 
* OUTPUT: fake_br_103 
* OUTPUT: fake_bl_104 
* OUTPUT: fake_br_104 
* OUTPUT: fake_bl_105 
* OUTPUT: fake_br_105 
* OUTPUT: fake_bl_106 
* OUTPUT: fake_br_106 
* OUTPUT: fake_bl_107 
* OUTPUT: fake_br_107 
* OUTPUT: fake_bl_108 
* OUTPUT: fake_br_108 
* OUTPUT: fake_bl_109 
* OUTPUT: fake_br_109 
* OUTPUT: fake_bl_110 
* OUTPUT: fake_br_110 
* OUTPUT: fake_bl_111 
* OUTPUT: fake_br_111 
* OUTPUT: fake_bl_112 
* OUTPUT: fake_br_112 
* OUTPUT: fake_bl_113 
* OUTPUT: fake_br_113 
* OUTPUT: fake_bl_114 
* OUTPUT: fake_br_114 
* OUTPUT: fake_bl_115 
* OUTPUT: fake_br_115 
* OUTPUT: fake_bl_116 
* OUTPUT: fake_br_116 
* OUTPUT: fake_bl_117 
* OUTPUT: fake_br_117 
* OUTPUT: fake_bl_118 
* OUTPUT: fake_br_118 
* OUTPUT: fake_bl_119 
* OUTPUT: fake_br_119 
* OUTPUT: fake_bl_120 
* OUTPUT: fake_br_120 
* OUTPUT: fake_bl_121 
* OUTPUT: fake_br_121 
* OUTPUT: fake_bl_122 
* OUTPUT: fake_br_122 
* OUTPUT: fake_bl_123 
* OUTPUT: fake_br_123 
* OUTPUT: fake_bl_124 
* OUTPUT: fake_br_124 
* OUTPUT: fake_bl_125 
* OUTPUT: fake_br_125 
* OUTPUT: fake_bl_126 
* OUTPUT: fake_br_126 
* OUTPUT: fake_bl_127 
* OUTPUT: fake_br_127 
* OUTPUT: fake_bl_128 
* OUTPUT: fake_br_128 
* INPUT : fake_wl 
* POWER : vdd 
* GROUND: gnd 
Xrca_top_0 fake_bl_0 vdd gnd fake_br_0 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_1 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_2 fake_bl_1 vdd gnd fake_br_1 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_3 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_4 fake_bl_2 vdd gnd fake_br_2 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_5 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_6 fake_bl_3 vdd gnd fake_br_3 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_7 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_8 fake_bl_4 vdd gnd fake_br_4 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_9 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_10 fake_bl_5 vdd gnd fake_br_5 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_11 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_12 fake_bl_6 vdd gnd fake_br_6 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_13 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_14 fake_bl_7 vdd gnd fake_br_7 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_15 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_16 fake_bl_8 vdd gnd fake_br_8 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_17 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_18 fake_bl_9 vdd gnd fake_br_9 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_19 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_20 fake_bl_10 vdd gnd fake_br_10 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_21 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_22 fake_bl_11 vdd gnd fake_br_11 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_23 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_24 fake_bl_12 vdd gnd fake_br_12 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_25 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_26 fake_bl_13 vdd gnd fake_br_13 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_27 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_28 fake_bl_14 vdd gnd fake_br_14 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_29 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_30 fake_bl_15 vdd gnd fake_br_15 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_31 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_32 fake_bl_16 vdd gnd fake_br_16 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_33 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_34 fake_bl_17 vdd gnd fake_br_17 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_35 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_36 fake_bl_18 vdd gnd fake_br_18 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_37 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_38 fake_bl_19 vdd gnd fake_br_19 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_39 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_40 fake_bl_20 vdd gnd fake_br_20 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_41 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_42 fake_bl_21 vdd gnd fake_br_21 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_43 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_44 fake_bl_22 vdd gnd fake_br_22 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_45 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_46 fake_bl_23 vdd gnd fake_br_23 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_47 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_48 fake_bl_24 vdd gnd fake_br_24 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_49 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_50 fake_bl_25 vdd gnd fake_br_25 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_51 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_52 fake_bl_26 vdd gnd fake_br_26 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_53 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_54 fake_bl_27 vdd gnd fake_br_27 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_55 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_56 fake_bl_28 vdd gnd fake_br_28 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_57 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_58 fake_bl_29 vdd gnd fake_br_29 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_59 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_60 fake_bl_30 vdd gnd fake_br_30 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_61 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_62 fake_bl_31 vdd gnd fake_br_31 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_63 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_64 fake_bl_32 vdd gnd fake_br_32 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_65 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_66 fake_bl_33 vdd gnd fake_br_33 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_67 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_68 fake_bl_34 vdd gnd fake_br_34 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_69 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_70 fake_bl_35 vdd gnd fake_br_35 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_71 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_72 fake_bl_36 vdd gnd fake_br_36 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_73 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_74 fake_bl_37 vdd gnd fake_br_37 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_75 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_76 fake_bl_38 vdd gnd fake_br_38 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_77 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_78 fake_bl_39 vdd gnd fake_br_39 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_79 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_80 fake_bl_40 vdd gnd fake_br_40 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_81 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_82 fake_bl_41 vdd gnd fake_br_41 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_83 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_84 fake_bl_42 vdd gnd fake_br_42 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_85 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_86 fake_bl_43 vdd gnd fake_br_43 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_87 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_88 fake_bl_44 vdd gnd fake_br_44 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_89 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_90 fake_bl_45 vdd gnd fake_br_45 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_91 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_92 fake_bl_46 vdd gnd fake_br_46 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_93 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_94 fake_bl_47 vdd gnd fake_br_47 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_95 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_96 fake_bl_48 vdd gnd fake_br_48 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_97 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_98 fake_bl_49 vdd gnd fake_br_49 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_99 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_100 fake_bl_50 vdd gnd fake_br_50 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_101 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_102 fake_bl_51 vdd gnd fake_br_51 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_103 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_104 fake_bl_52 vdd gnd fake_br_52 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_105 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_106 fake_bl_53 vdd gnd fake_br_53 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_107 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_108 fake_bl_54 vdd gnd fake_br_54 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_109 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_110 fake_bl_55 vdd gnd fake_br_55 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_111 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_112 fake_bl_56 vdd gnd fake_br_56 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_113 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_114 fake_bl_57 vdd gnd fake_br_57 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_115 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_116 fake_bl_58 vdd gnd fake_br_58 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_117 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_118 fake_bl_59 vdd gnd fake_br_59 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_119 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_120 fake_bl_60 vdd gnd fake_br_60 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_121 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_122 fake_bl_61 vdd gnd fake_br_61 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_123 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_124 fake_bl_62 vdd gnd fake_br_62 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_125 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_126 fake_bl_63 vdd gnd fake_br_63 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_127 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_128 fake_bl_64 vdd gnd fake_br_64 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_129 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_130 fake_bl_65 vdd gnd fake_br_65 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_131 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_132 fake_bl_66 vdd gnd fake_br_66 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_133 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_134 fake_bl_67 vdd gnd fake_br_67 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_135 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_136 fake_bl_68 vdd gnd fake_br_68 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_137 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_138 fake_bl_69 vdd gnd fake_br_69 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_139 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_140 fake_bl_70 vdd gnd fake_br_70 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_141 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_142 fake_bl_71 vdd gnd fake_br_71 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_143 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_144 fake_bl_72 vdd gnd fake_br_72 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_145 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_146 fake_bl_73 vdd gnd fake_br_73 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_147 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_148 fake_bl_74 vdd gnd fake_br_74 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_149 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_150 fake_bl_75 vdd gnd fake_br_75 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_151 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_152 fake_bl_76 vdd gnd fake_br_76 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_153 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_154 fake_bl_77 vdd gnd fake_br_77 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_155 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_156 fake_bl_78 vdd gnd fake_br_78 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_157 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_158 fake_bl_79 vdd gnd fake_br_79 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_159 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_160 fake_bl_80 vdd gnd fake_br_80 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_161 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_162 fake_bl_81 vdd gnd fake_br_81 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_163 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_164 fake_bl_82 vdd gnd fake_br_82 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_165 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_166 fake_bl_83 vdd gnd fake_br_83 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_167 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_168 fake_bl_84 vdd gnd fake_br_84 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_169 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_170 fake_bl_85 vdd gnd fake_br_85 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_171 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_172 fake_bl_86 vdd gnd fake_br_86 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_173 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_174 fake_bl_87 vdd gnd fake_br_87 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_175 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_176 fake_bl_88 vdd gnd fake_br_88 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_177 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_178 fake_bl_89 vdd gnd fake_br_89 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_179 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_180 fake_bl_90 vdd gnd fake_br_90 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_181 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_182 fake_bl_91 vdd gnd fake_br_91 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_183 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_184 fake_bl_92 vdd gnd fake_br_92 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_185 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_186 fake_bl_93 vdd gnd fake_br_93 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_187 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_188 fake_bl_94 vdd gnd fake_br_94 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_189 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_190 fake_bl_95 vdd gnd fake_br_95 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_191 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_192 fake_bl_96 vdd gnd fake_br_96 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_193 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_194 fake_bl_97 vdd gnd fake_br_97 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_195 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_196 fake_bl_98 vdd gnd fake_br_98 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_197 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_198 fake_bl_99 vdd gnd fake_br_99 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_199 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_200 fake_bl_100 vdd gnd fake_br_100 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_201 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_202 fake_bl_101 vdd gnd fake_br_101 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_203 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_204 fake_bl_102 vdd gnd fake_br_102 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_205 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_206 fake_bl_103 vdd gnd fake_br_103 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_207 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_208 fake_bl_104 vdd gnd fake_br_104 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_209 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_210 fake_bl_105 vdd gnd fake_br_105 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_211 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_212 fake_bl_106 vdd gnd fake_br_106 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_213 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_214 fake_bl_107 vdd gnd fake_br_107 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_215 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_216 fake_bl_108 vdd gnd fake_br_108 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_217 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_218 fake_bl_109 vdd gnd fake_br_109 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_219 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_220 fake_bl_110 vdd gnd fake_br_110 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_221 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_222 fake_bl_111 vdd gnd fake_br_111 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_223 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_224 fake_bl_112 vdd gnd fake_br_112 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_225 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_226 fake_bl_113 vdd gnd fake_br_113 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_227 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_228 fake_bl_114 vdd gnd fake_br_114 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_229 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_230 fake_bl_115 vdd gnd fake_br_115 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_231 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_232 fake_bl_116 vdd gnd fake_br_116 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_233 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_234 fake_bl_117 vdd gnd fake_br_117 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_235 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_236 fake_bl_118 vdd gnd fake_br_118 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_237 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_238 fake_bl_119 vdd gnd fake_br_119 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_239 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_240 fake_bl_120 vdd gnd fake_br_120 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_241 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_242 fake_bl_121 vdd gnd fake_br_121 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_243 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_244 fake_bl_122 vdd gnd fake_br_122 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_245 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_246 fake_bl_123 vdd gnd fake_br_123 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_247 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_248 fake_bl_124 vdd gnd fake_br_124 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_249 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_250 fake_bl_125 vdd gnd fake_br_125 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_251 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_252 fake_bl_126 vdd gnd fake_br_126 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_253 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_254 fake_bl_127 vdd gnd fake_br_127 sky130_fd_bd_sram__sram_sp_colend
Xrca_top_255 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_256 fake_bl_128 vdd gnd fake_br_128 sky130_fd_bd_sram__sram_sp_colend
.ENDS sky130_col_cap_array
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colenda_cent.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colenda_cent VPWR VPB VNB
.ends

.SUBCKT sky130_col_cap_array_0 fake_bl_0 fake_br_0 fake_bl_1 fake_br_1 fake_bl_2 fake_br_2 fake_bl_3 fake_br_3 fake_bl_4 fake_br_4 fake_bl_5 fake_br_5 fake_bl_6 fake_br_6 fake_bl_7 fake_br_7 fake_bl_8 fake_br_8 fake_bl_9 fake_br_9 fake_bl_10 fake_br_10 fake_bl_11 fake_br_11 fake_bl_12 fake_br_12 fake_bl_13 fake_br_13 fake_bl_14 fake_br_14 fake_bl_15 fake_br_15 fake_bl_16 fake_br_16 fake_bl_17 fake_br_17 fake_bl_18 fake_br_18 fake_bl_19 fake_br_19 fake_bl_20 fake_br_20 fake_bl_21 fake_br_21 fake_bl_22 fake_br_22 fake_bl_23 fake_br_23 fake_bl_24 fake_br_24 fake_bl_25 fake_br_25 fake_bl_26 fake_br_26 fake_bl_27 fake_br_27 fake_bl_28 fake_br_28 fake_bl_29 fake_br_29 fake_bl_30 fake_br_30 fake_bl_31 fake_br_31 fake_bl_32 fake_br_32 fake_bl_33 fake_br_33 fake_bl_34 fake_br_34 fake_bl_35 fake_br_35 fake_bl_36 fake_br_36 fake_bl_37 fake_br_37 fake_bl_38 fake_br_38 fake_bl_39 fake_br_39 fake_bl_40 fake_br_40 fake_bl_41 fake_br_41 fake_bl_42 fake_br_42 fake_bl_43 fake_br_43 fake_bl_44 fake_br_44 fake_bl_45 fake_br_45 fake_bl_46 fake_br_46 fake_bl_47 fake_br_47 fake_bl_48 fake_br_48 fake_bl_49 fake_br_49 fake_bl_50 fake_br_50 fake_bl_51 fake_br_51 fake_bl_52 fake_br_52 fake_bl_53 fake_br_53 fake_bl_54 fake_br_54 fake_bl_55 fake_br_55 fake_bl_56 fake_br_56 fake_bl_57 fake_br_57 fake_bl_58 fake_br_58 fake_bl_59 fake_br_59 fake_bl_60 fake_br_60 fake_bl_61 fake_br_61 fake_bl_62 fake_br_62 fake_bl_63 fake_br_63 fake_bl_64 fake_br_64 fake_bl_65 fake_br_65 fake_bl_66 fake_br_66 fake_bl_67 fake_br_67 fake_bl_68 fake_br_68 fake_bl_69 fake_br_69 fake_bl_70 fake_br_70 fake_bl_71 fake_br_71 fake_bl_72 fake_br_72 fake_bl_73 fake_br_73 fake_bl_74 fake_br_74 fake_bl_75 fake_br_75 fake_bl_76 fake_br_76 fake_bl_77 fake_br_77 fake_bl_78 fake_br_78 fake_bl_79 fake_br_79 fake_bl_80 fake_br_80 fake_bl_81 fake_br_81 fake_bl_82 fake_br_82 fake_bl_83 fake_br_83 fake_bl_84 fake_br_84 fake_bl_85 fake_br_85 fake_bl_86 fake_br_86 fake_bl_87 fake_br_87 fake_bl_88 fake_br_88 fake_bl_89 fake_br_89 fake_bl_90 fake_br_90 fake_bl_91 fake_br_91 fake_bl_92 fake_br_92 fake_bl_93 fake_br_93 fake_bl_94 fake_br_94 fake_bl_95 fake_br_95 fake_bl_96 fake_br_96 fake_bl_97 fake_br_97 fake_bl_98 fake_br_98 fake_bl_99 fake_br_99 fake_bl_100 fake_br_100 fake_bl_101 fake_br_101 fake_bl_102 fake_br_102 fake_bl_103 fake_br_103 fake_bl_104 fake_br_104 fake_bl_105 fake_br_105 fake_bl_106 fake_br_106 fake_bl_107 fake_br_107 fake_bl_108 fake_br_108 fake_bl_109 fake_br_109 fake_bl_110 fake_br_110 fake_bl_111 fake_br_111 fake_bl_112 fake_br_112 fake_bl_113 fake_br_113 fake_bl_114 fake_br_114 fake_bl_115 fake_br_115 fake_bl_116 fake_br_116 fake_bl_117 fake_br_117 fake_bl_118 fake_br_118 fake_bl_119 fake_br_119 fake_bl_120 fake_br_120 fake_bl_121 fake_br_121 fake_bl_122 fake_br_122 fake_bl_123 fake_br_123 fake_bl_124 fake_br_124 fake_bl_125 fake_br_125 fake_bl_126 fake_br_126 fake_bl_127 fake_br_127 fake_bl_128 fake_br_128 fake_wl vdd gnd
*.PININFO fake_bl_0:O fake_br_0:O fake_bl_1:O fake_br_1:O fake_bl_2:O fake_br_2:O fake_bl_3:O fake_br_3:O fake_bl_4:O fake_br_4:O fake_bl_5:O fake_br_5:O fake_bl_6:O fake_br_6:O fake_bl_7:O fake_br_7:O fake_bl_8:O fake_br_8:O fake_bl_9:O fake_br_9:O fake_bl_10:O fake_br_10:O fake_bl_11:O fake_br_11:O fake_bl_12:O fake_br_12:O fake_bl_13:O fake_br_13:O fake_bl_14:O fake_br_14:O fake_bl_15:O fake_br_15:O fake_bl_16:O fake_br_16:O fake_bl_17:O fake_br_17:O fake_bl_18:O fake_br_18:O fake_bl_19:O fake_br_19:O fake_bl_20:O fake_br_20:O fake_bl_21:O fake_br_21:O fake_bl_22:O fake_br_22:O fake_bl_23:O fake_br_23:O fake_bl_24:O fake_br_24:O fake_bl_25:O fake_br_25:O fake_bl_26:O fake_br_26:O fake_bl_27:O fake_br_27:O fake_bl_28:O fake_br_28:O fake_bl_29:O fake_br_29:O fake_bl_30:O fake_br_30:O fake_bl_31:O fake_br_31:O fake_bl_32:O fake_br_32:O fake_bl_33:O fake_br_33:O fake_bl_34:O fake_br_34:O fake_bl_35:O fake_br_35:O fake_bl_36:O fake_br_36:O fake_bl_37:O fake_br_37:O fake_bl_38:O fake_br_38:O fake_bl_39:O fake_br_39:O fake_bl_40:O fake_br_40:O fake_bl_41:O fake_br_41:O fake_bl_42:O fake_br_42:O fake_bl_43:O fake_br_43:O fake_bl_44:O fake_br_44:O fake_bl_45:O fake_br_45:O fake_bl_46:O fake_br_46:O fake_bl_47:O fake_br_47:O fake_bl_48:O fake_br_48:O fake_bl_49:O fake_br_49:O fake_bl_50:O fake_br_50:O fake_bl_51:O fake_br_51:O fake_bl_52:O fake_br_52:O fake_bl_53:O fake_br_53:O fake_bl_54:O fake_br_54:O fake_bl_55:O fake_br_55:O fake_bl_56:O fake_br_56:O fake_bl_57:O fake_br_57:O fake_bl_58:O fake_br_58:O fake_bl_59:O fake_br_59:O fake_bl_60:O fake_br_60:O fake_bl_61:O fake_br_61:O fake_bl_62:O fake_br_62:O fake_bl_63:O fake_br_63:O fake_bl_64:O fake_br_64:O fake_bl_65:O fake_br_65:O fake_bl_66:O fake_br_66:O fake_bl_67:O fake_br_67:O fake_bl_68:O fake_br_68:O fake_bl_69:O fake_br_69:O fake_bl_70:O fake_br_70:O fake_bl_71:O fake_br_71:O fake_bl_72:O fake_br_72:O fake_bl_73:O fake_br_73:O fake_bl_74:O fake_br_74:O fake_bl_75:O fake_br_75:O fake_bl_76:O fake_br_76:O fake_bl_77:O fake_br_77:O fake_bl_78:O fake_br_78:O fake_bl_79:O fake_br_79:O fake_bl_80:O fake_br_80:O fake_bl_81:O fake_br_81:O fake_bl_82:O fake_br_82:O fake_bl_83:O fake_br_83:O fake_bl_84:O fake_br_84:O fake_bl_85:O fake_br_85:O fake_bl_86:O fake_br_86:O fake_bl_87:O fake_br_87:O fake_bl_88:O fake_br_88:O fake_bl_89:O fake_br_89:O fake_bl_90:O fake_br_90:O fake_bl_91:O fake_br_91:O fake_bl_92:O fake_br_92:O fake_bl_93:O fake_br_93:O fake_bl_94:O fake_br_94:O fake_bl_95:O fake_br_95:O fake_bl_96:O fake_br_96:O fake_bl_97:O fake_br_97:O fake_bl_98:O fake_br_98:O fake_bl_99:O fake_br_99:O fake_bl_100:O fake_br_100:O fake_bl_101:O fake_br_101:O fake_bl_102:O fake_br_102:O fake_bl_103:O fake_br_103:O fake_bl_104:O fake_br_104:O fake_bl_105:O fake_br_105:O fake_bl_106:O fake_br_106:O fake_bl_107:O fake_br_107:O fake_bl_108:O fake_br_108:O fake_bl_109:O fake_br_109:O fake_bl_110:O fake_br_110:O fake_bl_111:O fake_br_111:O fake_bl_112:O fake_br_112:O fake_bl_113:O fake_br_113:O fake_bl_114:O fake_br_114:O fake_bl_115:O fake_br_115:O fake_bl_116:O fake_br_116:O fake_bl_117:O fake_br_117:O fake_bl_118:O fake_br_118:O fake_bl_119:O fake_br_119:O fake_bl_120:O fake_br_120:O fake_bl_121:O fake_br_121:O fake_bl_122:O fake_br_122:O fake_bl_123:O fake_br_123:O fake_bl_124:O fake_br_124:O fake_bl_125:O fake_br_125:O fake_bl_126:O fake_br_126:O fake_bl_127:O fake_br_127:O fake_bl_128:O fake_br_128:O fake_wl:I vdd:B gnd:B
* OUTPUT: fake_bl_0 
* OUTPUT: fake_br_0 
* OUTPUT: fake_bl_1 
* OUTPUT: fake_br_1 
* OUTPUT: fake_bl_2 
* OUTPUT: fake_br_2 
* OUTPUT: fake_bl_3 
* OUTPUT: fake_br_3 
* OUTPUT: fake_bl_4 
* OUTPUT: fake_br_4 
* OUTPUT: fake_bl_5 
* OUTPUT: fake_br_5 
* OUTPUT: fake_bl_6 
* OUTPUT: fake_br_6 
* OUTPUT: fake_bl_7 
* OUTPUT: fake_br_7 
* OUTPUT: fake_bl_8 
* OUTPUT: fake_br_8 
* OUTPUT: fake_bl_9 
* OUTPUT: fake_br_9 
* OUTPUT: fake_bl_10 
* OUTPUT: fake_br_10 
* OUTPUT: fake_bl_11 
* OUTPUT: fake_br_11 
* OUTPUT: fake_bl_12 
* OUTPUT: fake_br_12 
* OUTPUT: fake_bl_13 
* OUTPUT: fake_br_13 
* OUTPUT: fake_bl_14 
* OUTPUT: fake_br_14 
* OUTPUT: fake_bl_15 
* OUTPUT: fake_br_15 
* OUTPUT: fake_bl_16 
* OUTPUT: fake_br_16 
* OUTPUT: fake_bl_17 
* OUTPUT: fake_br_17 
* OUTPUT: fake_bl_18 
* OUTPUT: fake_br_18 
* OUTPUT: fake_bl_19 
* OUTPUT: fake_br_19 
* OUTPUT: fake_bl_20 
* OUTPUT: fake_br_20 
* OUTPUT: fake_bl_21 
* OUTPUT: fake_br_21 
* OUTPUT: fake_bl_22 
* OUTPUT: fake_br_22 
* OUTPUT: fake_bl_23 
* OUTPUT: fake_br_23 
* OUTPUT: fake_bl_24 
* OUTPUT: fake_br_24 
* OUTPUT: fake_bl_25 
* OUTPUT: fake_br_25 
* OUTPUT: fake_bl_26 
* OUTPUT: fake_br_26 
* OUTPUT: fake_bl_27 
* OUTPUT: fake_br_27 
* OUTPUT: fake_bl_28 
* OUTPUT: fake_br_28 
* OUTPUT: fake_bl_29 
* OUTPUT: fake_br_29 
* OUTPUT: fake_bl_30 
* OUTPUT: fake_br_30 
* OUTPUT: fake_bl_31 
* OUTPUT: fake_br_31 
* OUTPUT: fake_bl_32 
* OUTPUT: fake_br_32 
* OUTPUT: fake_bl_33 
* OUTPUT: fake_br_33 
* OUTPUT: fake_bl_34 
* OUTPUT: fake_br_34 
* OUTPUT: fake_bl_35 
* OUTPUT: fake_br_35 
* OUTPUT: fake_bl_36 
* OUTPUT: fake_br_36 
* OUTPUT: fake_bl_37 
* OUTPUT: fake_br_37 
* OUTPUT: fake_bl_38 
* OUTPUT: fake_br_38 
* OUTPUT: fake_bl_39 
* OUTPUT: fake_br_39 
* OUTPUT: fake_bl_40 
* OUTPUT: fake_br_40 
* OUTPUT: fake_bl_41 
* OUTPUT: fake_br_41 
* OUTPUT: fake_bl_42 
* OUTPUT: fake_br_42 
* OUTPUT: fake_bl_43 
* OUTPUT: fake_br_43 
* OUTPUT: fake_bl_44 
* OUTPUT: fake_br_44 
* OUTPUT: fake_bl_45 
* OUTPUT: fake_br_45 
* OUTPUT: fake_bl_46 
* OUTPUT: fake_br_46 
* OUTPUT: fake_bl_47 
* OUTPUT: fake_br_47 
* OUTPUT: fake_bl_48 
* OUTPUT: fake_br_48 
* OUTPUT: fake_bl_49 
* OUTPUT: fake_br_49 
* OUTPUT: fake_bl_50 
* OUTPUT: fake_br_50 
* OUTPUT: fake_bl_51 
* OUTPUT: fake_br_51 
* OUTPUT: fake_bl_52 
* OUTPUT: fake_br_52 
* OUTPUT: fake_bl_53 
* OUTPUT: fake_br_53 
* OUTPUT: fake_bl_54 
* OUTPUT: fake_br_54 
* OUTPUT: fake_bl_55 
* OUTPUT: fake_br_55 
* OUTPUT: fake_bl_56 
* OUTPUT: fake_br_56 
* OUTPUT: fake_bl_57 
* OUTPUT: fake_br_57 
* OUTPUT: fake_bl_58 
* OUTPUT: fake_br_58 
* OUTPUT: fake_bl_59 
* OUTPUT: fake_br_59 
* OUTPUT: fake_bl_60 
* OUTPUT: fake_br_60 
* OUTPUT: fake_bl_61 
* OUTPUT: fake_br_61 
* OUTPUT: fake_bl_62 
* OUTPUT: fake_br_62 
* OUTPUT: fake_bl_63 
* OUTPUT: fake_br_63 
* OUTPUT: fake_bl_64 
* OUTPUT: fake_br_64 
* OUTPUT: fake_bl_65 
* OUTPUT: fake_br_65 
* OUTPUT: fake_bl_66 
* OUTPUT: fake_br_66 
* OUTPUT: fake_bl_67 
* OUTPUT: fake_br_67 
* OUTPUT: fake_bl_68 
* OUTPUT: fake_br_68 
* OUTPUT: fake_bl_69 
* OUTPUT: fake_br_69 
* OUTPUT: fake_bl_70 
* OUTPUT: fake_br_70 
* OUTPUT: fake_bl_71 
* OUTPUT: fake_br_71 
* OUTPUT: fake_bl_72 
* OUTPUT: fake_br_72 
* OUTPUT: fake_bl_73 
* OUTPUT: fake_br_73 
* OUTPUT: fake_bl_74 
* OUTPUT: fake_br_74 
* OUTPUT: fake_bl_75 
* OUTPUT: fake_br_75 
* OUTPUT: fake_bl_76 
* OUTPUT: fake_br_76 
* OUTPUT: fake_bl_77 
* OUTPUT: fake_br_77 
* OUTPUT: fake_bl_78 
* OUTPUT: fake_br_78 
* OUTPUT: fake_bl_79 
* OUTPUT: fake_br_79 
* OUTPUT: fake_bl_80 
* OUTPUT: fake_br_80 
* OUTPUT: fake_bl_81 
* OUTPUT: fake_br_81 
* OUTPUT: fake_bl_82 
* OUTPUT: fake_br_82 
* OUTPUT: fake_bl_83 
* OUTPUT: fake_br_83 
* OUTPUT: fake_bl_84 
* OUTPUT: fake_br_84 
* OUTPUT: fake_bl_85 
* OUTPUT: fake_br_85 
* OUTPUT: fake_bl_86 
* OUTPUT: fake_br_86 
* OUTPUT: fake_bl_87 
* OUTPUT: fake_br_87 
* OUTPUT: fake_bl_88 
* OUTPUT: fake_br_88 
* OUTPUT: fake_bl_89 
* OUTPUT: fake_br_89 
* OUTPUT: fake_bl_90 
* OUTPUT: fake_br_90 
* OUTPUT: fake_bl_91 
* OUTPUT: fake_br_91 
* OUTPUT: fake_bl_92 
* OUTPUT: fake_br_92 
* OUTPUT: fake_bl_93 
* OUTPUT: fake_br_93 
* OUTPUT: fake_bl_94 
* OUTPUT: fake_br_94 
* OUTPUT: fake_bl_95 
* OUTPUT: fake_br_95 
* OUTPUT: fake_bl_96 
* OUTPUT: fake_br_96 
* OUTPUT: fake_bl_97 
* OUTPUT: fake_br_97 
* OUTPUT: fake_bl_98 
* OUTPUT: fake_br_98 
* OUTPUT: fake_bl_99 
* OUTPUT: fake_br_99 
* OUTPUT: fake_bl_100 
* OUTPUT: fake_br_100 
* OUTPUT: fake_bl_101 
* OUTPUT: fake_br_101 
* OUTPUT: fake_bl_102 
* OUTPUT: fake_br_102 
* OUTPUT: fake_bl_103 
* OUTPUT: fake_br_103 
* OUTPUT: fake_bl_104 
* OUTPUT: fake_br_104 
* OUTPUT: fake_bl_105 
* OUTPUT: fake_br_105 
* OUTPUT: fake_bl_106 
* OUTPUT: fake_br_106 
* OUTPUT: fake_bl_107 
* OUTPUT: fake_br_107 
* OUTPUT: fake_bl_108 
* OUTPUT: fake_br_108 
* OUTPUT: fake_bl_109 
* OUTPUT: fake_br_109 
* OUTPUT: fake_bl_110 
* OUTPUT: fake_br_110 
* OUTPUT: fake_bl_111 
* OUTPUT: fake_br_111 
* OUTPUT: fake_bl_112 
* OUTPUT: fake_br_112 
* OUTPUT: fake_bl_113 
* OUTPUT: fake_br_113 
* OUTPUT: fake_bl_114 
* OUTPUT: fake_br_114 
* OUTPUT: fake_bl_115 
* OUTPUT: fake_br_115 
* OUTPUT: fake_bl_116 
* OUTPUT: fake_br_116 
* OUTPUT: fake_bl_117 
* OUTPUT: fake_br_117 
* OUTPUT: fake_bl_118 
* OUTPUT: fake_br_118 
* OUTPUT: fake_bl_119 
* OUTPUT: fake_br_119 
* OUTPUT: fake_bl_120 
* OUTPUT: fake_br_120 
* OUTPUT: fake_bl_121 
* OUTPUT: fake_br_121 
* OUTPUT: fake_bl_122 
* OUTPUT: fake_br_122 
* OUTPUT: fake_bl_123 
* OUTPUT: fake_br_123 
* OUTPUT: fake_bl_124 
* OUTPUT: fake_br_124 
* OUTPUT: fake_bl_125 
* OUTPUT: fake_br_125 
* OUTPUT: fake_bl_126 
* OUTPUT: fake_br_126 
* OUTPUT: fake_bl_127 
* OUTPUT: fake_br_127 
* OUTPUT: fake_bl_128 
* OUTPUT: fake_br_128 
* INPUT : fake_wl 
* POWER : vdd 
* GROUND: gnd 
Xrca_bottom_0 fake_bl_0 vdd gnd fake_br_0 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_1 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_2 fake_bl_1 vdd gnd fake_br_1 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_3 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_4 fake_bl_2 vdd gnd fake_br_2 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_5 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_6 fake_bl_3 vdd gnd fake_br_3 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_7 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_8 fake_bl_4 vdd gnd fake_br_4 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_9 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_10 fake_bl_5 vdd gnd fake_br_5 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_11 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_12 fake_bl_6 vdd gnd fake_br_6 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_13 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_14 fake_bl_7 vdd gnd fake_br_7 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_15 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_16 fake_bl_8 vdd gnd fake_br_8 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_17 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_18 fake_bl_9 vdd gnd fake_br_9 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_19 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_20 fake_bl_10 vdd gnd fake_br_10 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_21 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_22 fake_bl_11 vdd gnd fake_br_11 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_23 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_24 fake_bl_12 vdd gnd fake_br_12 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_25 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_26 fake_bl_13 vdd gnd fake_br_13 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_27 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_28 fake_bl_14 vdd gnd fake_br_14 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_29 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_30 fake_bl_15 vdd gnd fake_br_15 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_31 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_32 fake_bl_16 vdd gnd fake_br_16 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_33 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_34 fake_bl_17 vdd gnd fake_br_17 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_35 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_36 fake_bl_18 vdd gnd fake_br_18 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_37 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_38 fake_bl_19 vdd gnd fake_br_19 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_39 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_40 fake_bl_20 vdd gnd fake_br_20 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_41 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_42 fake_bl_21 vdd gnd fake_br_21 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_43 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_44 fake_bl_22 vdd gnd fake_br_22 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_45 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_46 fake_bl_23 vdd gnd fake_br_23 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_47 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_48 fake_bl_24 vdd gnd fake_br_24 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_49 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_50 fake_bl_25 vdd gnd fake_br_25 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_51 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_52 fake_bl_26 vdd gnd fake_br_26 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_53 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_54 fake_bl_27 vdd gnd fake_br_27 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_55 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_56 fake_bl_28 vdd gnd fake_br_28 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_57 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_58 fake_bl_29 vdd gnd fake_br_29 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_59 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_60 fake_bl_30 vdd gnd fake_br_30 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_61 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_62 fake_bl_31 vdd gnd fake_br_31 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_63 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_64 fake_bl_32 vdd gnd fake_br_32 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_65 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_66 fake_bl_33 vdd gnd fake_br_33 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_67 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_68 fake_bl_34 vdd gnd fake_br_34 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_69 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_70 fake_bl_35 vdd gnd fake_br_35 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_71 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_72 fake_bl_36 vdd gnd fake_br_36 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_73 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_74 fake_bl_37 vdd gnd fake_br_37 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_75 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_76 fake_bl_38 vdd gnd fake_br_38 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_77 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_78 fake_bl_39 vdd gnd fake_br_39 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_79 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_80 fake_bl_40 vdd gnd fake_br_40 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_81 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_82 fake_bl_41 vdd gnd fake_br_41 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_83 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_84 fake_bl_42 vdd gnd fake_br_42 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_85 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_86 fake_bl_43 vdd gnd fake_br_43 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_87 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_88 fake_bl_44 vdd gnd fake_br_44 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_89 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_90 fake_bl_45 vdd gnd fake_br_45 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_91 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_92 fake_bl_46 vdd gnd fake_br_46 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_93 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_94 fake_bl_47 vdd gnd fake_br_47 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_95 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_96 fake_bl_48 vdd gnd fake_br_48 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_97 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_98 fake_bl_49 vdd gnd fake_br_49 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_99 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_100 fake_bl_50 vdd gnd fake_br_50 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_101 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_102 fake_bl_51 vdd gnd fake_br_51 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_103 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_104 fake_bl_52 vdd gnd fake_br_52 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_105 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_106 fake_bl_53 vdd gnd fake_br_53 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_107 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_108 fake_bl_54 vdd gnd fake_br_54 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_109 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_110 fake_bl_55 vdd gnd fake_br_55 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_111 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_112 fake_bl_56 vdd gnd fake_br_56 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_113 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_114 fake_bl_57 vdd gnd fake_br_57 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_115 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_116 fake_bl_58 vdd gnd fake_br_58 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_117 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_118 fake_bl_59 vdd gnd fake_br_59 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_119 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_120 fake_bl_60 vdd gnd fake_br_60 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_121 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_122 fake_bl_61 vdd gnd fake_br_61 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_123 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_124 fake_bl_62 vdd gnd fake_br_62 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_125 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_126 fake_bl_63 vdd gnd fake_br_63 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_127 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_128 fake_bl_64 vdd gnd fake_br_64 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_129 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_130 fake_bl_65 vdd gnd fake_br_65 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_131 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_132 fake_bl_66 vdd gnd fake_br_66 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_133 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_134 fake_bl_67 vdd gnd fake_br_67 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_135 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_136 fake_bl_68 vdd gnd fake_br_68 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_137 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_138 fake_bl_69 vdd gnd fake_br_69 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_139 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_140 fake_bl_70 vdd gnd fake_br_70 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_141 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_142 fake_bl_71 vdd gnd fake_br_71 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_143 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_144 fake_bl_72 vdd gnd fake_br_72 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_145 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_146 fake_bl_73 vdd gnd fake_br_73 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_147 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_148 fake_bl_74 vdd gnd fake_br_74 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_149 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_150 fake_bl_75 vdd gnd fake_br_75 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_151 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_152 fake_bl_76 vdd gnd fake_br_76 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_153 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_154 fake_bl_77 vdd gnd fake_br_77 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_155 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_156 fake_bl_78 vdd gnd fake_br_78 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_157 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_158 fake_bl_79 vdd gnd fake_br_79 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_159 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_160 fake_bl_80 vdd gnd fake_br_80 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_161 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_162 fake_bl_81 vdd gnd fake_br_81 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_163 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_164 fake_bl_82 vdd gnd fake_br_82 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_165 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_166 fake_bl_83 vdd gnd fake_br_83 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_167 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_168 fake_bl_84 vdd gnd fake_br_84 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_169 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_170 fake_bl_85 vdd gnd fake_br_85 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_171 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_172 fake_bl_86 vdd gnd fake_br_86 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_173 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_174 fake_bl_87 vdd gnd fake_br_87 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_175 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_176 fake_bl_88 vdd gnd fake_br_88 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_177 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_178 fake_bl_89 vdd gnd fake_br_89 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_179 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_180 fake_bl_90 vdd gnd fake_br_90 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_181 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_182 fake_bl_91 vdd gnd fake_br_91 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_183 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_184 fake_bl_92 vdd gnd fake_br_92 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_185 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_186 fake_bl_93 vdd gnd fake_br_93 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_187 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_188 fake_bl_94 vdd gnd fake_br_94 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_189 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_190 fake_bl_95 vdd gnd fake_br_95 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_191 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_192 fake_bl_96 vdd gnd fake_br_96 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_193 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_194 fake_bl_97 vdd gnd fake_br_97 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_195 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_196 fake_bl_98 vdd gnd fake_br_98 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_197 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_198 fake_bl_99 vdd gnd fake_br_99 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_199 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_200 fake_bl_100 vdd gnd fake_br_100 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_201 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_202 fake_bl_101 vdd gnd fake_br_101 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_203 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_204 fake_bl_102 vdd gnd fake_br_102 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_205 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_206 fake_bl_103 vdd gnd fake_br_103 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_207 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_208 fake_bl_104 vdd gnd fake_br_104 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_209 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_210 fake_bl_105 vdd gnd fake_br_105 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_211 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_212 fake_bl_106 vdd gnd fake_br_106 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_213 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_214 fake_bl_107 vdd gnd fake_br_107 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_215 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_216 fake_bl_108 vdd gnd fake_br_108 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_217 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_218 fake_bl_109 vdd gnd fake_br_109 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_219 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_220 fake_bl_110 vdd gnd fake_br_110 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_221 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_222 fake_bl_111 vdd gnd fake_br_111 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_223 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_224 fake_bl_112 vdd gnd fake_br_112 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_225 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_226 fake_bl_113 vdd gnd fake_br_113 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_227 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_228 fake_bl_114 vdd gnd fake_br_114 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_229 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_230 fake_bl_115 vdd gnd fake_br_115 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_231 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_232 fake_bl_116 vdd gnd fake_br_116 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_233 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_234 fake_bl_117 vdd gnd fake_br_117 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_235 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_236 fake_bl_118 vdd gnd fake_br_118 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_237 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_238 fake_bl_119 vdd gnd fake_br_119 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_239 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_240 fake_bl_120 vdd gnd fake_br_120 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_241 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_242 fake_bl_121 vdd gnd fake_br_121 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_243 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_244 fake_bl_122 vdd gnd fake_br_122 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_245 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_246 fake_bl_123 vdd gnd fake_br_123 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_247 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_248 fake_bl_124 vdd gnd fake_br_124 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_249 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_250 fake_bl_125 vdd gnd fake_br_125 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_251 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_252 fake_bl_126 vdd gnd fake_br_126 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_253 vdd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_254 fake_bl_127 vdd gnd fake_br_127 sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_255 gnd vdd gnd sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_256 fake_bl_128 vdd gnd fake_br_128 sky130_fd_bd_sram__sram_sp_colenda
.ENDS sky130_col_cap_array_0
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_corner.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_corner VPWR VPB VNB
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_cornera.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_cornera VNB VPWR VPB
.ends
* NGSPICE file created from sky130_fd_bd_sram__openram_sp_rowend_replica.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_rowend_replica VPWR WL
.ends
* NGSPICE file created from sky130_fd_bd_sram__openram_sp_rowenda_replica.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_rowenda_replica VPWR WL
.ends

.SUBCKT sky130_row_cap_array wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 wl_0_129 wl_0_130 wl_0_131 vdd gnd
*.PININFO wl_0_0:O wl_0_1:O wl_0_2:O wl_0_3:O wl_0_4:O wl_0_5:O wl_0_6:O wl_0_7:O wl_0_8:O wl_0_9:O wl_0_10:O wl_0_11:O wl_0_12:O wl_0_13:O wl_0_14:O wl_0_15:O wl_0_16:O wl_0_17:O wl_0_18:O wl_0_19:O wl_0_20:O wl_0_21:O wl_0_22:O wl_0_23:O wl_0_24:O wl_0_25:O wl_0_26:O wl_0_27:O wl_0_28:O wl_0_29:O wl_0_30:O wl_0_31:O wl_0_32:O wl_0_33:O wl_0_34:O wl_0_35:O wl_0_36:O wl_0_37:O wl_0_38:O wl_0_39:O wl_0_40:O wl_0_41:O wl_0_42:O wl_0_43:O wl_0_44:O wl_0_45:O wl_0_46:O wl_0_47:O wl_0_48:O wl_0_49:O wl_0_50:O wl_0_51:O wl_0_52:O wl_0_53:O wl_0_54:O wl_0_55:O wl_0_56:O wl_0_57:O wl_0_58:O wl_0_59:O wl_0_60:O wl_0_61:O wl_0_62:O wl_0_63:O wl_0_64:O wl_0_65:O wl_0_66:O wl_0_67:O wl_0_68:O wl_0_69:O wl_0_70:O wl_0_71:O wl_0_72:O wl_0_73:O wl_0_74:O wl_0_75:O wl_0_76:O wl_0_77:O wl_0_78:O wl_0_79:O wl_0_80:O wl_0_81:O wl_0_82:O wl_0_83:O wl_0_84:O wl_0_85:O wl_0_86:O wl_0_87:O wl_0_88:O wl_0_89:O wl_0_90:O wl_0_91:O wl_0_92:O wl_0_93:O wl_0_94:O wl_0_95:O wl_0_96:O wl_0_97:O wl_0_98:O wl_0_99:O wl_0_100:O wl_0_101:O wl_0_102:O wl_0_103:O wl_0_104:O wl_0_105:O wl_0_106:O wl_0_107:O wl_0_108:O wl_0_109:O wl_0_110:O wl_0_111:O wl_0_112:O wl_0_113:O wl_0_114:O wl_0_115:O wl_0_116:O wl_0_117:O wl_0_118:O wl_0_119:O wl_0_120:O wl_0_121:O wl_0_122:O wl_0_123:O wl_0_124:O wl_0_125:O wl_0_126:O wl_0_127:O wl_0_128:O wl_0_129:O wl_0_130:O wl_0_131:O vdd:B gnd:B
* OUTPUT: wl_0_0 
* OUTPUT: wl_0_1 
* OUTPUT: wl_0_2 
* OUTPUT: wl_0_3 
* OUTPUT: wl_0_4 
* OUTPUT: wl_0_5 
* OUTPUT: wl_0_6 
* OUTPUT: wl_0_7 
* OUTPUT: wl_0_8 
* OUTPUT: wl_0_9 
* OUTPUT: wl_0_10 
* OUTPUT: wl_0_11 
* OUTPUT: wl_0_12 
* OUTPUT: wl_0_13 
* OUTPUT: wl_0_14 
* OUTPUT: wl_0_15 
* OUTPUT: wl_0_16 
* OUTPUT: wl_0_17 
* OUTPUT: wl_0_18 
* OUTPUT: wl_0_19 
* OUTPUT: wl_0_20 
* OUTPUT: wl_0_21 
* OUTPUT: wl_0_22 
* OUTPUT: wl_0_23 
* OUTPUT: wl_0_24 
* OUTPUT: wl_0_25 
* OUTPUT: wl_0_26 
* OUTPUT: wl_0_27 
* OUTPUT: wl_0_28 
* OUTPUT: wl_0_29 
* OUTPUT: wl_0_30 
* OUTPUT: wl_0_31 
* OUTPUT: wl_0_32 
* OUTPUT: wl_0_33 
* OUTPUT: wl_0_34 
* OUTPUT: wl_0_35 
* OUTPUT: wl_0_36 
* OUTPUT: wl_0_37 
* OUTPUT: wl_0_38 
* OUTPUT: wl_0_39 
* OUTPUT: wl_0_40 
* OUTPUT: wl_0_41 
* OUTPUT: wl_0_42 
* OUTPUT: wl_0_43 
* OUTPUT: wl_0_44 
* OUTPUT: wl_0_45 
* OUTPUT: wl_0_46 
* OUTPUT: wl_0_47 
* OUTPUT: wl_0_48 
* OUTPUT: wl_0_49 
* OUTPUT: wl_0_50 
* OUTPUT: wl_0_51 
* OUTPUT: wl_0_52 
* OUTPUT: wl_0_53 
* OUTPUT: wl_0_54 
* OUTPUT: wl_0_55 
* OUTPUT: wl_0_56 
* OUTPUT: wl_0_57 
* OUTPUT: wl_0_58 
* OUTPUT: wl_0_59 
* OUTPUT: wl_0_60 
* OUTPUT: wl_0_61 
* OUTPUT: wl_0_62 
* OUTPUT: wl_0_63 
* OUTPUT: wl_0_64 
* OUTPUT: wl_0_65 
* OUTPUT: wl_0_66 
* OUTPUT: wl_0_67 
* OUTPUT: wl_0_68 
* OUTPUT: wl_0_69 
* OUTPUT: wl_0_70 
* OUTPUT: wl_0_71 
* OUTPUT: wl_0_72 
* OUTPUT: wl_0_73 
* OUTPUT: wl_0_74 
* OUTPUT: wl_0_75 
* OUTPUT: wl_0_76 
* OUTPUT: wl_0_77 
* OUTPUT: wl_0_78 
* OUTPUT: wl_0_79 
* OUTPUT: wl_0_80 
* OUTPUT: wl_0_81 
* OUTPUT: wl_0_82 
* OUTPUT: wl_0_83 
* OUTPUT: wl_0_84 
* OUTPUT: wl_0_85 
* OUTPUT: wl_0_86 
* OUTPUT: wl_0_87 
* OUTPUT: wl_0_88 
* OUTPUT: wl_0_89 
* OUTPUT: wl_0_90 
* OUTPUT: wl_0_91 
* OUTPUT: wl_0_92 
* OUTPUT: wl_0_93 
* OUTPUT: wl_0_94 
* OUTPUT: wl_0_95 
* OUTPUT: wl_0_96 
* OUTPUT: wl_0_97 
* OUTPUT: wl_0_98 
* OUTPUT: wl_0_99 
* OUTPUT: wl_0_100 
* OUTPUT: wl_0_101 
* OUTPUT: wl_0_102 
* OUTPUT: wl_0_103 
* OUTPUT: wl_0_104 
* OUTPUT: wl_0_105 
* OUTPUT: wl_0_106 
* OUTPUT: wl_0_107 
* OUTPUT: wl_0_108 
* OUTPUT: wl_0_109 
* OUTPUT: wl_0_110 
* OUTPUT: wl_0_111 
* OUTPUT: wl_0_112 
* OUTPUT: wl_0_113 
* OUTPUT: wl_0_114 
* OUTPUT: wl_0_115 
* OUTPUT: wl_0_116 
* OUTPUT: wl_0_117 
* OUTPUT: wl_0_118 
* OUTPUT: wl_0_119 
* OUTPUT: wl_0_120 
* OUTPUT: wl_0_121 
* OUTPUT: wl_0_122 
* OUTPUT: wl_0_123 
* OUTPUT: wl_0_124 
* OUTPUT: wl_0_125 
* OUTPUT: wl_0_126 
* OUTPUT: wl_0_127 
* OUTPUT: wl_0_128 
* OUTPUT: wl_0_129 
* OUTPUT: wl_0_130 
* OUTPUT: wl_0_131 
* POWER : vdd 
* GROUND: gnd 
Xrca_0 vdd gnd vdd sky130_fd_bd_sram__sram_sp_cornera
Xrca_1 wl_0_0 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_2 wl_0_1 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_3 wl_0_2 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_4 wl_0_3 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_5 wl_0_4 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_6 wl_0_5 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_7 wl_0_6 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_8 wl_0_7 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_9 wl_0_8 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_10 wl_0_9 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_11 wl_0_10 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_12 wl_0_11 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_13 wl_0_12 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_14 wl_0_13 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_15 wl_0_14 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_16 wl_0_15 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_17 wl_0_16 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_18 wl_0_17 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_19 wl_0_18 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_20 wl_0_19 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_21 wl_0_20 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_22 wl_0_21 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_23 wl_0_22 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_24 wl_0_23 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_25 wl_0_24 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_26 wl_0_25 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_27 wl_0_26 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_28 wl_0_27 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_29 wl_0_28 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_30 wl_0_29 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_31 wl_0_30 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_32 wl_0_31 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_33 wl_0_32 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_34 wl_0_33 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_35 wl_0_34 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_36 wl_0_35 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_37 wl_0_36 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_38 wl_0_37 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_39 wl_0_38 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_40 wl_0_39 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_41 wl_0_40 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_42 wl_0_41 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_43 wl_0_42 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_44 wl_0_43 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_45 wl_0_44 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_46 wl_0_45 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_47 wl_0_46 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_48 wl_0_47 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_49 wl_0_48 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_50 wl_0_49 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_51 wl_0_50 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_52 wl_0_51 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_53 wl_0_52 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_54 wl_0_53 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_55 wl_0_54 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_56 wl_0_55 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_57 wl_0_56 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_58 wl_0_57 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_59 wl_0_58 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_60 wl_0_59 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_61 wl_0_60 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_62 wl_0_61 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_63 wl_0_62 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_64 wl_0_63 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_65 wl_0_64 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_66 wl_0_65 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_67 wl_0_66 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_68 wl_0_67 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_69 wl_0_68 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_70 wl_0_69 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_71 wl_0_70 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_72 wl_0_71 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_73 wl_0_72 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_74 wl_0_73 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_75 wl_0_74 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_76 wl_0_75 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_77 wl_0_76 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_78 wl_0_77 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_79 wl_0_78 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_80 wl_0_79 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_81 wl_0_80 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_82 wl_0_81 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_83 wl_0_82 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_84 wl_0_83 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_85 wl_0_84 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_86 wl_0_85 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_87 wl_0_86 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_88 wl_0_87 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_89 wl_0_88 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_90 wl_0_89 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_91 wl_0_90 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_92 wl_0_91 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_93 wl_0_92 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_94 wl_0_93 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_95 wl_0_94 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_96 wl_0_95 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_97 wl_0_96 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_98 wl_0_97 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_99 wl_0_98 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_100 wl_0_99 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_101 wl_0_100 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_102 wl_0_101 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_103 wl_0_102 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_104 wl_0_103 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_105 wl_0_104 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_106 wl_0_105 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_107 wl_0_106 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_108 wl_0_107 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_109 wl_0_108 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_110 wl_0_109 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_111 wl_0_110 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_112 wl_0_111 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_113 wl_0_112 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_114 wl_0_113 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_115 wl_0_114 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_116 wl_0_115 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_117 wl_0_116 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_118 wl_0_117 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_119 wl_0_118 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_120 wl_0_119 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_121 wl_0_120 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_122 wl_0_121 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_123 wl_0_122 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_124 wl_0_123 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_125 wl_0_124 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_126 wl_0_125 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_127 wl_0_126 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_128 wl_0_127 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_129 wl_0_128 vdd sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_130 wl_0_129 vdd sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_131 vdd gnd vdd sky130_fd_bd_sram__sram_sp_corner
.ENDS sky130_row_cap_array
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_cornerb.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_cornerb VPWR VPB VNB
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_rowend.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_rowend VPWR WL
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_rowenda.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_rowenda VPWR WL
.ends

.SUBCKT sky130_row_cap_array_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 wl_0_129 wl_0_130 wl_0_131 vdd gnd
*.PININFO wl_0_0:O wl_0_1:O wl_0_2:O wl_0_3:O wl_0_4:O wl_0_5:O wl_0_6:O wl_0_7:O wl_0_8:O wl_0_9:O wl_0_10:O wl_0_11:O wl_0_12:O wl_0_13:O wl_0_14:O wl_0_15:O wl_0_16:O wl_0_17:O wl_0_18:O wl_0_19:O wl_0_20:O wl_0_21:O wl_0_22:O wl_0_23:O wl_0_24:O wl_0_25:O wl_0_26:O wl_0_27:O wl_0_28:O wl_0_29:O wl_0_30:O wl_0_31:O wl_0_32:O wl_0_33:O wl_0_34:O wl_0_35:O wl_0_36:O wl_0_37:O wl_0_38:O wl_0_39:O wl_0_40:O wl_0_41:O wl_0_42:O wl_0_43:O wl_0_44:O wl_0_45:O wl_0_46:O wl_0_47:O wl_0_48:O wl_0_49:O wl_0_50:O wl_0_51:O wl_0_52:O wl_0_53:O wl_0_54:O wl_0_55:O wl_0_56:O wl_0_57:O wl_0_58:O wl_0_59:O wl_0_60:O wl_0_61:O wl_0_62:O wl_0_63:O wl_0_64:O wl_0_65:O wl_0_66:O wl_0_67:O wl_0_68:O wl_0_69:O wl_0_70:O wl_0_71:O wl_0_72:O wl_0_73:O wl_0_74:O wl_0_75:O wl_0_76:O wl_0_77:O wl_0_78:O wl_0_79:O wl_0_80:O wl_0_81:O wl_0_82:O wl_0_83:O wl_0_84:O wl_0_85:O wl_0_86:O wl_0_87:O wl_0_88:O wl_0_89:O wl_0_90:O wl_0_91:O wl_0_92:O wl_0_93:O wl_0_94:O wl_0_95:O wl_0_96:O wl_0_97:O wl_0_98:O wl_0_99:O wl_0_100:O wl_0_101:O wl_0_102:O wl_0_103:O wl_0_104:O wl_0_105:O wl_0_106:O wl_0_107:O wl_0_108:O wl_0_109:O wl_0_110:O wl_0_111:O wl_0_112:O wl_0_113:O wl_0_114:O wl_0_115:O wl_0_116:O wl_0_117:O wl_0_118:O wl_0_119:O wl_0_120:O wl_0_121:O wl_0_122:O wl_0_123:O wl_0_124:O wl_0_125:O wl_0_126:O wl_0_127:O wl_0_128:O wl_0_129:O wl_0_130:O wl_0_131:O vdd:B gnd:B
* OUTPUT: wl_0_0 
* OUTPUT: wl_0_1 
* OUTPUT: wl_0_2 
* OUTPUT: wl_0_3 
* OUTPUT: wl_0_4 
* OUTPUT: wl_0_5 
* OUTPUT: wl_0_6 
* OUTPUT: wl_0_7 
* OUTPUT: wl_0_8 
* OUTPUT: wl_0_9 
* OUTPUT: wl_0_10 
* OUTPUT: wl_0_11 
* OUTPUT: wl_0_12 
* OUTPUT: wl_0_13 
* OUTPUT: wl_0_14 
* OUTPUT: wl_0_15 
* OUTPUT: wl_0_16 
* OUTPUT: wl_0_17 
* OUTPUT: wl_0_18 
* OUTPUT: wl_0_19 
* OUTPUT: wl_0_20 
* OUTPUT: wl_0_21 
* OUTPUT: wl_0_22 
* OUTPUT: wl_0_23 
* OUTPUT: wl_0_24 
* OUTPUT: wl_0_25 
* OUTPUT: wl_0_26 
* OUTPUT: wl_0_27 
* OUTPUT: wl_0_28 
* OUTPUT: wl_0_29 
* OUTPUT: wl_0_30 
* OUTPUT: wl_0_31 
* OUTPUT: wl_0_32 
* OUTPUT: wl_0_33 
* OUTPUT: wl_0_34 
* OUTPUT: wl_0_35 
* OUTPUT: wl_0_36 
* OUTPUT: wl_0_37 
* OUTPUT: wl_0_38 
* OUTPUT: wl_0_39 
* OUTPUT: wl_0_40 
* OUTPUT: wl_0_41 
* OUTPUT: wl_0_42 
* OUTPUT: wl_0_43 
* OUTPUT: wl_0_44 
* OUTPUT: wl_0_45 
* OUTPUT: wl_0_46 
* OUTPUT: wl_0_47 
* OUTPUT: wl_0_48 
* OUTPUT: wl_0_49 
* OUTPUT: wl_0_50 
* OUTPUT: wl_0_51 
* OUTPUT: wl_0_52 
* OUTPUT: wl_0_53 
* OUTPUT: wl_0_54 
* OUTPUT: wl_0_55 
* OUTPUT: wl_0_56 
* OUTPUT: wl_0_57 
* OUTPUT: wl_0_58 
* OUTPUT: wl_0_59 
* OUTPUT: wl_0_60 
* OUTPUT: wl_0_61 
* OUTPUT: wl_0_62 
* OUTPUT: wl_0_63 
* OUTPUT: wl_0_64 
* OUTPUT: wl_0_65 
* OUTPUT: wl_0_66 
* OUTPUT: wl_0_67 
* OUTPUT: wl_0_68 
* OUTPUT: wl_0_69 
* OUTPUT: wl_0_70 
* OUTPUT: wl_0_71 
* OUTPUT: wl_0_72 
* OUTPUT: wl_0_73 
* OUTPUT: wl_0_74 
* OUTPUT: wl_0_75 
* OUTPUT: wl_0_76 
* OUTPUT: wl_0_77 
* OUTPUT: wl_0_78 
* OUTPUT: wl_0_79 
* OUTPUT: wl_0_80 
* OUTPUT: wl_0_81 
* OUTPUT: wl_0_82 
* OUTPUT: wl_0_83 
* OUTPUT: wl_0_84 
* OUTPUT: wl_0_85 
* OUTPUT: wl_0_86 
* OUTPUT: wl_0_87 
* OUTPUT: wl_0_88 
* OUTPUT: wl_0_89 
* OUTPUT: wl_0_90 
* OUTPUT: wl_0_91 
* OUTPUT: wl_0_92 
* OUTPUT: wl_0_93 
* OUTPUT: wl_0_94 
* OUTPUT: wl_0_95 
* OUTPUT: wl_0_96 
* OUTPUT: wl_0_97 
* OUTPUT: wl_0_98 
* OUTPUT: wl_0_99 
* OUTPUT: wl_0_100 
* OUTPUT: wl_0_101 
* OUTPUT: wl_0_102 
* OUTPUT: wl_0_103 
* OUTPUT: wl_0_104 
* OUTPUT: wl_0_105 
* OUTPUT: wl_0_106 
* OUTPUT: wl_0_107 
* OUTPUT: wl_0_108 
* OUTPUT: wl_0_109 
* OUTPUT: wl_0_110 
* OUTPUT: wl_0_111 
* OUTPUT: wl_0_112 
* OUTPUT: wl_0_113 
* OUTPUT: wl_0_114 
* OUTPUT: wl_0_115 
* OUTPUT: wl_0_116 
* OUTPUT: wl_0_117 
* OUTPUT: wl_0_118 
* OUTPUT: wl_0_119 
* OUTPUT: wl_0_120 
* OUTPUT: wl_0_121 
* OUTPUT: wl_0_122 
* OUTPUT: wl_0_123 
* OUTPUT: wl_0_124 
* OUTPUT: wl_0_125 
* OUTPUT: wl_0_126 
* OUTPUT: wl_0_127 
* OUTPUT: wl_0_128 
* OUTPUT: wl_0_129 
* OUTPUT: wl_0_130 
* OUTPUT: wl_0_131 
* POWER : vdd 
* GROUND: gnd 
Xrca_0 vdd gnd vdd sky130_fd_bd_sram__sram_sp_cornera
Xrca_1 wl_0_0 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_2 wl_0_1 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_3 wl_0_2 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_4 wl_0_3 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_5 wl_0_4 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_6 wl_0_5 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_7 wl_0_6 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_8 wl_0_7 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_9 wl_0_8 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_10 wl_0_9 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_11 wl_0_10 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_12 wl_0_11 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_13 wl_0_12 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_14 wl_0_13 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_15 wl_0_14 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_16 wl_0_15 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_17 wl_0_16 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_18 wl_0_17 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_19 wl_0_18 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_20 wl_0_19 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_21 wl_0_20 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_22 wl_0_21 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_23 wl_0_22 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_24 wl_0_23 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_25 wl_0_24 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_26 wl_0_25 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_27 wl_0_26 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_28 wl_0_27 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_29 wl_0_28 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_30 wl_0_29 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_31 wl_0_30 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_32 wl_0_31 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_33 wl_0_32 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_34 wl_0_33 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_35 wl_0_34 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_36 wl_0_35 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_37 wl_0_36 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_38 wl_0_37 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_39 wl_0_38 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_40 wl_0_39 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_41 wl_0_40 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_42 wl_0_41 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_43 wl_0_42 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_44 wl_0_43 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_45 wl_0_44 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_46 wl_0_45 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_47 wl_0_46 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_48 wl_0_47 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_49 wl_0_48 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_50 wl_0_49 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_51 wl_0_50 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_52 wl_0_51 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_53 wl_0_52 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_54 wl_0_53 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_55 wl_0_54 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_56 wl_0_55 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_57 wl_0_56 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_58 wl_0_57 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_59 wl_0_58 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_60 wl_0_59 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_61 wl_0_60 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_62 wl_0_61 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_63 wl_0_62 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_64 wl_0_63 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_65 wl_0_64 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_66 wl_0_65 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_67 wl_0_66 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_68 wl_0_67 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_69 wl_0_68 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_70 wl_0_69 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_71 wl_0_70 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_72 wl_0_71 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_73 wl_0_72 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_74 wl_0_73 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_75 wl_0_74 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_76 wl_0_75 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_77 wl_0_76 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_78 wl_0_77 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_79 wl_0_78 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_80 wl_0_79 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_81 wl_0_80 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_82 wl_0_81 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_83 wl_0_82 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_84 wl_0_83 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_85 wl_0_84 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_86 wl_0_85 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_87 wl_0_86 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_88 wl_0_87 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_89 wl_0_88 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_90 wl_0_89 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_91 wl_0_90 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_92 wl_0_91 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_93 wl_0_92 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_94 wl_0_93 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_95 wl_0_94 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_96 wl_0_95 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_97 wl_0_96 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_98 wl_0_97 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_99 wl_0_98 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_100 wl_0_99 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_101 wl_0_100 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_102 wl_0_101 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_103 wl_0_102 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_104 wl_0_103 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_105 wl_0_104 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_106 wl_0_105 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_107 wl_0_106 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_108 wl_0_107 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_109 wl_0_108 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_110 wl_0_109 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_111 wl_0_110 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_112 wl_0_111 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_113 wl_0_112 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_114 wl_0_113 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_115 wl_0_114 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_116 wl_0_115 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_117 wl_0_116 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_118 wl_0_117 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_119 wl_0_118 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_120 wl_0_119 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_121 wl_0_120 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_122 wl_0_121 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_123 wl_0_122 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_124 wl_0_123 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_125 wl_0_124 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_126 wl_0_125 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_127 wl_0_126 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_128 wl_0_127 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_129 wl_0_128 vdd sky130_fd_bd_sram__sram_sp_rowenda
Xrca_130 wl_0_129 vdd sky130_fd_bd_sram__sram_sp_rowend
Xrca_131 vdd gnd vdd sky130_fd_bd_sram__sram_sp_cornerb
.ENDS sky130_row_cap_array_0

.SUBCKT sky130_replica_bitcell_array rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 vdd gnd vpb vnb
*.PININFO rbl_bl_0_0:B rbl_br_0_0:B bl_0_0:B br_0_0:B bl_0_1:B br_0_1:B bl_0_2:B br_0_2:B bl_0_3:B br_0_3:B bl_0_4:B br_0_4:B bl_0_5:B br_0_5:B bl_0_6:B br_0_6:B bl_0_7:B br_0_7:B bl_0_8:B br_0_8:B bl_0_9:B br_0_9:B bl_0_10:B br_0_10:B bl_0_11:B br_0_11:B bl_0_12:B br_0_12:B bl_0_13:B br_0_13:B bl_0_14:B br_0_14:B bl_0_15:B br_0_15:B bl_0_16:B br_0_16:B bl_0_17:B br_0_17:B bl_0_18:B br_0_18:B bl_0_19:B br_0_19:B bl_0_20:B br_0_20:B bl_0_21:B br_0_21:B bl_0_22:B br_0_22:B bl_0_23:B br_0_23:B bl_0_24:B br_0_24:B bl_0_25:B br_0_25:B bl_0_26:B br_0_26:B bl_0_27:B br_0_27:B bl_0_28:B br_0_28:B bl_0_29:B br_0_29:B bl_0_30:B br_0_30:B bl_0_31:B br_0_31:B bl_0_32:B br_0_32:B bl_0_33:B br_0_33:B bl_0_34:B br_0_34:B bl_0_35:B br_0_35:B bl_0_36:B br_0_36:B bl_0_37:B br_0_37:B bl_0_38:B br_0_38:B bl_0_39:B br_0_39:B bl_0_40:B br_0_40:B bl_0_41:B br_0_41:B bl_0_42:B br_0_42:B bl_0_43:B br_0_43:B bl_0_44:B br_0_44:B bl_0_45:B br_0_45:B bl_0_46:B br_0_46:B bl_0_47:B br_0_47:B bl_0_48:B br_0_48:B bl_0_49:B br_0_49:B bl_0_50:B br_0_50:B bl_0_51:B br_0_51:B bl_0_52:B br_0_52:B bl_0_53:B br_0_53:B bl_0_54:B br_0_54:B bl_0_55:B br_0_55:B bl_0_56:B br_0_56:B bl_0_57:B br_0_57:B bl_0_58:B br_0_58:B bl_0_59:B br_0_59:B bl_0_60:B br_0_60:B bl_0_61:B br_0_61:B bl_0_62:B br_0_62:B bl_0_63:B br_0_63:B bl_0_64:B br_0_64:B bl_0_65:B br_0_65:B bl_0_66:B br_0_66:B bl_0_67:B br_0_67:B bl_0_68:B br_0_68:B bl_0_69:B br_0_69:B bl_0_70:B br_0_70:B bl_0_71:B br_0_71:B bl_0_72:B br_0_72:B bl_0_73:B br_0_73:B bl_0_74:B br_0_74:B bl_0_75:B br_0_75:B bl_0_76:B br_0_76:B bl_0_77:B br_0_77:B bl_0_78:B br_0_78:B bl_0_79:B br_0_79:B bl_0_80:B br_0_80:B bl_0_81:B br_0_81:B bl_0_82:B br_0_82:B bl_0_83:B br_0_83:B bl_0_84:B br_0_84:B bl_0_85:B br_0_85:B bl_0_86:B br_0_86:B bl_0_87:B br_0_87:B bl_0_88:B br_0_88:B bl_0_89:B br_0_89:B bl_0_90:B br_0_90:B bl_0_91:B br_0_91:B bl_0_92:B br_0_92:B bl_0_93:B br_0_93:B bl_0_94:B br_0_94:B bl_0_95:B br_0_95:B bl_0_96:B br_0_96:B bl_0_97:B br_0_97:B bl_0_98:B br_0_98:B bl_0_99:B br_0_99:B bl_0_100:B br_0_100:B bl_0_101:B br_0_101:B bl_0_102:B br_0_102:B bl_0_103:B br_0_103:B bl_0_104:B br_0_104:B bl_0_105:B br_0_105:B bl_0_106:B br_0_106:B bl_0_107:B br_0_107:B bl_0_108:B br_0_108:B bl_0_109:B br_0_109:B bl_0_110:B br_0_110:B bl_0_111:B br_0_111:B bl_0_112:B br_0_112:B bl_0_113:B br_0_113:B bl_0_114:B br_0_114:B bl_0_115:B br_0_115:B bl_0_116:B br_0_116:B bl_0_117:B br_0_117:B bl_0_118:B br_0_118:B bl_0_119:B br_0_119:B bl_0_120:B br_0_120:B bl_0_121:B br_0_121:B bl_0_122:B br_0_122:B bl_0_123:B br_0_123:B bl_0_124:B br_0_124:B bl_0_125:B br_0_125:B bl_0_126:B br_0_126:B bl_0_127:B br_0_127:B bl_0_128:B br_0_128:B rbl_wl_0_0:I wl_0_0:I wl_0_1:I wl_0_2:I wl_0_3:I wl_0_4:I wl_0_5:I wl_0_6:I wl_0_7:I wl_0_8:I wl_0_9:I wl_0_10:I wl_0_11:I wl_0_12:I wl_0_13:I wl_0_14:I wl_0_15:I wl_0_16:I wl_0_17:I wl_0_18:I wl_0_19:I wl_0_20:I wl_0_21:I wl_0_22:I wl_0_23:I wl_0_24:I wl_0_25:I wl_0_26:I wl_0_27:I wl_0_28:I wl_0_29:I wl_0_30:I wl_0_31:I wl_0_32:I wl_0_33:I wl_0_34:I wl_0_35:I wl_0_36:I wl_0_37:I wl_0_38:I wl_0_39:I wl_0_40:I wl_0_41:I wl_0_42:I wl_0_43:I wl_0_44:I wl_0_45:I wl_0_46:I wl_0_47:I wl_0_48:I wl_0_49:I wl_0_50:I wl_0_51:I wl_0_52:I wl_0_53:I wl_0_54:I wl_0_55:I wl_0_56:I wl_0_57:I wl_0_58:I wl_0_59:I wl_0_60:I wl_0_61:I wl_0_62:I wl_0_63:I wl_0_64:I wl_0_65:I wl_0_66:I wl_0_67:I wl_0_68:I wl_0_69:I wl_0_70:I wl_0_71:I wl_0_72:I wl_0_73:I wl_0_74:I wl_0_75:I wl_0_76:I wl_0_77:I wl_0_78:I wl_0_79:I wl_0_80:I wl_0_81:I wl_0_82:I wl_0_83:I wl_0_84:I wl_0_85:I wl_0_86:I wl_0_87:I wl_0_88:I wl_0_89:I wl_0_90:I wl_0_91:I wl_0_92:I wl_0_93:I wl_0_94:I wl_0_95:I wl_0_96:I wl_0_97:I wl_0_98:I wl_0_99:I wl_0_100:I wl_0_101:I wl_0_102:I wl_0_103:I wl_0_104:I wl_0_105:I wl_0_106:I wl_0_107:I wl_0_108:I wl_0_109:I wl_0_110:I wl_0_111:I wl_0_112:I wl_0_113:I wl_0_114:I wl_0_115:I wl_0_116:I wl_0_117:I wl_0_118:I wl_0_119:I wl_0_120:I wl_0_121:I wl_0_122:I wl_0_123:I wl_0_124:I wl_0_125:I wl_0_126:I wl_0_127:I wl_0_128:I vdd:B gnd:B vpb:B vnb:B
* INOUT : rbl_bl_0_0 
* INOUT : rbl_br_0_0 
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INPUT : rbl_wl_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* INPUT : wl_0_67 
* INPUT : wl_0_68 
* INPUT : wl_0_69 
* INPUT : wl_0_70 
* INPUT : wl_0_71 
* INPUT : wl_0_72 
* INPUT : wl_0_73 
* INPUT : wl_0_74 
* INPUT : wl_0_75 
* INPUT : wl_0_76 
* INPUT : wl_0_77 
* INPUT : wl_0_78 
* INPUT : wl_0_79 
* INPUT : wl_0_80 
* INPUT : wl_0_81 
* INPUT : wl_0_82 
* INPUT : wl_0_83 
* INPUT : wl_0_84 
* INPUT : wl_0_85 
* INPUT : wl_0_86 
* INPUT : wl_0_87 
* INPUT : wl_0_88 
* INPUT : wl_0_89 
* INPUT : wl_0_90 
* INPUT : wl_0_91 
* INPUT : wl_0_92 
* INPUT : wl_0_93 
* INPUT : wl_0_94 
* INPUT : wl_0_95 
* INPUT : wl_0_96 
* INPUT : wl_0_97 
* INPUT : wl_0_98 
* INPUT : wl_0_99 
* INPUT : wl_0_100 
* INPUT : wl_0_101 
* INPUT : wl_0_102 
* INPUT : wl_0_103 
* INPUT : wl_0_104 
* INPUT : wl_0_105 
* INPUT : wl_0_106 
* INPUT : wl_0_107 
* INPUT : wl_0_108 
* INPUT : wl_0_109 
* INPUT : wl_0_110 
* INPUT : wl_0_111 
* INPUT : wl_0_112 
* INPUT : wl_0_113 
* INPUT : wl_0_114 
* INPUT : wl_0_115 
* INPUT : wl_0_116 
* INPUT : wl_0_117 
* INPUT : wl_0_118 
* INPUT : wl_0_119 
* INPUT : wl_0_120 
* INPUT : wl_0_121 
* INPUT : wl_0_122 
* INPUT : wl_0_123 
* INPUT : wl_0_124 
* INPUT : wl_0_125 
* INPUT : wl_0_126 
* INPUT : wl_0_127 
* INPUT : wl_0_128 
* POWER : vdd 
* GROUND: gnd 
* BIAS  : vpb 
* BIAS  : vnb 
* rbl: None left_rbl: None right_rbl: None
Xbitcell_array bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 vdd gnd sky130_bitcell_array
Xreplica_col_0 rbl_bl_0_0 rbl_br_0_0 gnd rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 gnd vdd gnd sky130_replica_column
Xdummy_row_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 rbl_wl_0_0 vdd gnd sky130_dummy_array
Xdummy_row_bot bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 gnd vdd gnd sky130_col_cap_array_0
Xdummy_row_top bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 gnd vdd gnd sky130_col_cap_array
Xdummy_col_left gnd rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 gnd vdd gnd sky130_row_cap_array
Xdummy_col_right gnd rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 gnd vdd gnd sky130_row_cap_array_0
.ENDS sky130_replica_bitcell_array
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* NGSPICE file created from sky130_fd_bd_sram__openram_sp_nand2_dec.ext - technology: EFS8A


* Top level circuit sky130_fd_bd_sram__openram_sp_nand2_dec
.subckt sky130_fd_bd_sram__openram_sp_nand2_dec A B Z VDD GND

X1001 Z B VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1002 VDD A Z VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1000 Z A a_n722_276# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1003 a_n722_276# B GND GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
.ends


* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u

.SUBCKT pinv_dec A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS pinv_dec

.SUBCKT and2_dec A B Z vdd gnd
*.PININFO A:I B:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand2_dec_nand A B zb_int vdd gnd sky130_fd_bd_sram__openram_sp_nand2_dec
Xpand2_dec_inv zb_int Z vdd gnd pinv_dec
.ENDS and2_dec
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* NGSPICE file created from sky130_fd_bd_sram__openram_sp_nand3_dec.ext - technology: EFS8A


* Top level circuit sky130_fd_bd_sram__openram_sp_nand3_dec
.subckt sky130_fd_bd_sram__openram_sp_nand3_dec A B C Z VDD GND

X1001 Z A a_n346_328# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1002 a_n346_256# C GND GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1003 a_n346_328# B a_n346_256# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1000 Z B VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1004 Z A VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1005 Z C VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
.ends


.SUBCKT and3_dec A B C Z vdd gnd
*.PININFO A:I B:I C:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand3_dec_nand A B C zb_int vdd gnd sky130_fd_bd_sram__openram_sp_nand3_dec
Xpand3_dec_inv zb_int Z vdd gnd pinv_dec
.ENDS and3_dec

.SUBCKT hierarchical_predecode2x4 in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
*.PININFO in_0:I in_1:I out_0:O out_1:O out_2:O out_3:O vdd:B gnd:B
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_dec
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_dec
XXpre2x4_and_0 inbar_0 inbar_1 out_0 vdd gnd and2_dec
XXpre2x4_and_1 in_0 inbar_1 out_1 vdd gnd and2_dec
XXpre2x4_and_2 inbar_0 in_1 out_2 vdd gnd and2_dec
XXpre2x4_and_3 in_0 in_1 out_3 vdd gnd and2_dec
.ENDS hierarchical_predecode2x4

.SUBCKT hierarchical_predecode3x8 in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
*.PININFO in_0:I in_1:I in_2:I out_0:O out_1:O out_2:O out_3:O out_4:O out_5:O out_6:O out_7:O vdd:B gnd:B
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_dec
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_dec
Xpre_inv_2 in_2 inbar_2 vdd gnd pinv_dec
XXpre3x8_and_0 inbar_0 inbar_1 inbar_2 out_0 vdd gnd and3_dec
XXpre3x8_and_1 in_0 inbar_1 inbar_2 out_1 vdd gnd and3_dec
XXpre3x8_and_2 inbar_0 in_1 inbar_2 out_2 vdd gnd and3_dec
XXpre3x8_and_3 in_0 in_1 inbar_2 out_3 vdd gnd and3_dec
XXpre3x8_and_4 inbar_0 inbar_1 in_2 out_4 vdd gnd and3_dec
XXpre3x8_and_5 in_0 inbar_1 in_2 out_5 vdd gnd and3_dec
XXpre3x8_and_6 inbar_0 in_1 in_2 out_6 vdd gnd and3_dec
XXpre3x8_and_7 in_0 in_1 in_2 out_7 vdd gnd and3_dec
.ENDS hierarchical_predecode3x8
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* NGSPICE file created from sky130_fd_bd_sram__openram_sp_nand4_dec.ext - technology: EFS8A

.subckt sky130_fd_bd_sram__openram_sp_nand4_dec A B C D Z VDD GND
X1000 Z A a_406_334# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1004 a_406_190# D GND GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1005 a_406_262# C a_406_190# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1007 a_406_334# B a_406_262# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1001 Z A VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1002 VDD C Z VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1003 VDD D Z VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1006 Z B VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
.ends


.SUBCKT and4_dec A B C D Z vdd gnd
*.PININFO A:I B:I C:I D:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* INPUT : C 
* INPUT : D 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand4_dec_nand A B C D zb_int vdd gnd sky130_fd_bd_sram__openram_sp_nand4_dec
Xpand4_dec_inv zb_int Z vdd gnd pinv_dec
.ENDS and4_dec

.SUBCKT hierarchical_predecode4x16 in_0 in_1 in_2 in_3 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 out_8 out_9 out_10 out_11 out_12 out_13 out_14 out_15 vdd gnd
*.PININFO in_0:I in_1:I in_2:I in_3:I out_0:O out_1:O out_2:O out_3:O out_4:O out_5:O out_6:O out_7:O out_8:O out_9:O out_10:O out_11:O out_12:O out_13:O out_14:O out_15:O vdd:B gnd:B
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* OUTPUT: out_8 
* OUTPUT: out_9 
* OUTPUT: out_10 
* OUTPUT: out_11 
* OUTPUT: out_12 
* OUTPUT: out_13 
* OUTPUT: out_14 
* OUTPUT: out_15 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_dec
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_dec
Xpre_inv_2 in_2 inbar_2 vdd gnd pinv_dec
Xpre_inv_3 in_3 inbar_3 vdd gnd pinv_dec
XXpre4x16_and_0 inbar_0 inbar_1 inbar_2 inbar_3 out_0 vdd gnd and4_dec
XXpre4x16_and_1 in_0 inbar_1 inbar_2 inbar_3 out_1 vdd gnd and4_dec
XXpre4x16_and_2 inbar_0 in_1 inbar_2 inbar_3 out_2 vdd gnd and4_dec
XXpre4x16_and_3 in_0 in_1 inbar_2 inbar_3 out_3 vdd gnd and4_dec
XXpre4x16_and_4 inbar_0 inbar_1 in_2 inbar_3 out_4 vdd gnd and4_dec
XXpre4x16_and_5 in_0 inbar_1 in_2 inbar_3 out_5 vdd gnd and4_dec
XXpre4x16_and_6 inbar_0 in_1 in_2 inbar_3 out_6 vdd gnd and4_dec
XXpre4x16_and_7 in_0 in_1 in_2 inbar_3 out_7 vdd gnd and4_dec
XXpre4x16_and_8 inbar_0 inbar_1 inbar_2 in_3 out_8 vdd gnd and4_dec
XXpre4x16_and_9 in_0 inbar_1 inbar_2 in_3 out_9 vdd gnd and4_dec
XXpre4x16_and_10 inbar_0 in_1 inbar_2 in_3 out_10 vdd gnd and4_dec
XXpre4x16_and_11 in_0 in_1 inbar_2 in_3 out_11 vdd gnd and4_dec
XXpre4x16_and_12 inbar_0 inbar_1 in_2 in_3 out_12 vdd gnd and4_dec
XXpre4x16_and_13 in_0 inbar_1 in_2 in_3 out_13 vdd gnd and4_dec
XXpre4x16_and_14 inbar_0 in_1 in_2 in_3 out_14 vdd gnd and4_dec
XXpre4x16_and_15 in_0 in_1 in_2 in_3 out_15 vdd gnd and4_dec
.ENDS hierarchical_predecode4x16

.SUBCKT hierarchical_decoder addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 addr_7 decode_0 decode_1 decode_2 decode_3 decode_4 decode_5 decode_6 decode_7 decode_8 decode_9 decode_10 decode_11 decode_12 decode_13 decode_14 decode_15 decode_16 decode_17 decode_18 decode_19 decode_20 decode_21 decode_22 decode_23 decode_24 decode_25 decode_26 decode_27 decode_28 decode_29 decode_30 decode_31 decode_32 decode_33 decode_34 decode_35 decode_36 decode_37 decode_38 decode_39 decode_40 decode_41 decode_42 decode_43 decode_44 decode_45 decode_46 decode_47 decode_48 decode_49 decode_50 decode_51 decode_52 decode_53 decode_54 decode_55 decode_56 decode_57 decode_58 decode_59 decode_60 decode_61 decode_62 decode_63 decode_64 decode_65 decode_66 decode_67 decode_68 decode_69 decode_70 decode_71 decode_72 decode_73 decode_74 decode_75 decode_76 decode_77 decode_78 decode_79 decode_80 decode_81 decode_82 decode_83 decode_84 decode_85 decode_86 decode_87 decode_88 decode_89 decode_90 decode_91 decode_92 decode_93 decode_94 decode_95 decode_96 decode_97 decode_98 decode_99 decode_100 decode_101 decode_102 decode_103 decode_104 decode_105 decode_106 decode_107 decode_108 decode_109 decode_110 decode_111 decode_112 decode_113 decode_114 decode_115 decode_116 decode_117 decode_118 decode_119 decode_120 decode_121 decode_122 decode_123 decode_124 decode_125 decode_126 decode_127 decode_128 vdd gnd
*.PININFO addr_0:I addr_1:I addr_2:I addr_3:I addr_4:I addr_5:I addr_6:I addr_7:I decode_0:O decode_1:O decode_2:O decode_3:O decode_4:O decode_5:O decode_6:O decode_7:O decode_8:O decode_9:O decode_10:O decode_11:O decode_12:O decode_13:O decode_14:O decode_15:O decode_16:O decode_17:O decode_18:O decode_19:O decode_20:O decode_21:O decode_22:O decode_23:O decode_24:O decode_25:O decode_26:O decode_27:O decode_28:O decode_29:O decode_30:O decode_31:O decode_32:O decode_33:O decode_34:O decode_35:O decode_36:O decode_37:O decode_38:O decode_39:O decode_40:O decode_41:O decode_42:O decode_43:O decode_44:O decode_45:O decode_46:O decode_47:O decode_48:O decode_49:O decode_50:O decode_51:O decode_52:O decode_53:O decode_54:O decode_55:O decode_56:O decode_57:O decode_58:O decode_59:O decode_60:O decode_61:O decode_62:O decode_63:O decode_64:O decode_65:O decode_66:O decode_67:O decode_68:O decode_69:O decode_70:O decode_71:O decode_72:O decode_73:O decode_74:O decode_75:O decode_76:O decode_77:O decode_78:O decode_79:O decode_80:O decode_81:O decode_82:O decode_83:O decode_84:O decode_85:O decode_86:O decode_87:O decode_88:O decode_89:O decode_90:O decode_91:O decode_92:O decode_93:O decode_94:O decode_95:O decode_96:O decode_97:O decode_98:O decode_99:O decode_100:O decode_101:O decode_102:O decode_103:O decode_104:O decode_105:O decode_106:O decode_107:O decode_108:O decode_109:O decode_110:O decode_111:O decode_112:O decode_113:O decode_114:O decode_115:O decode_116:O decode_117:O decode_118:O decode_119:O decode_120:O decode_121:O decode_122:O decode_123:O decode_124:O decode_125:O decode_126:O decode_127:O decode_128:O vdd:B gnd:B
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* INPUT : addr_7 
* OUTPUT: decode_0 
* OUTPUT: decode_1 
* OUTPUT: decode_2 
* OUTPUT: decode_3 
* OUTPUT: decode_4 
* OUTPUT: decode_5 
* OUTPUT: decode_6 
* OUTPUT: decode_7 
* OUTPUT: decode_8 
* OUTPUT: decode_9 
* OUTPUT: decode_10 
* OUTPUT: decode_11 
* OUTPUT: decode_12 
* OUTPUT: decode_13 
* OUTPUT: decode_14 
* OUTPUT: decode_15 
* OUTPUT: decode_16 
* OUTPUT: decode_17 
* OUTPUT: decode_18 
* OUTPUT: decode_19 
* OUTPUT: decode_20 
* OUTPUT: decode_21 
* OUTPUT: decode_22 
* OUTPUT: decode_23 
* OUTPUT: decode_24 
* OUTPUT: decode_25 
* OUTPUT: decode_26 
* OUTPUT: decode_27 
* OUTPUT: decode_28 
* OUTPUT: decode_29 
* OUTPUT: decode_30 
* OUTPUT: decode_31 
* OUTPUT: decode_32 
* OUTPUT: decode_33 
* OUTPUT: decode_34 
* OUTPUT: decode_35 
* OUTPUT: decode_36 
* OUTPUT: decode_37 
* OUTPUT: decode_38 
* OUTPUT: decode_39 
* OUTPUT: decode_40 
* OUTPUT: decode_41 
* OUTPUT: decode_42 
* OUTPUT: decode_43 
* OUTPUT: decode_44 
* OUTPUT: decode_45 
* OUTPUT: decode_46 
* OUTPUT: decode_47 
* OUTPUT: decode_48 
* OUTPUT: decode_49 
* OUTPUT: decode_50 
* OUTPUT: decode_51 
* OUTPUT: decode_52 
* OUTPUT: decode_53 
* OUTPUT: decode_54 
* OUTPUT: decode_55 
* OUTPUT: decode_56 
* OUTPUT: decode_57 
* OUTPUT: decode_58 
* OUTPUT: decode_59 
* OUTPUT: decode_60 
* OUTPUT: decode_61 
* OUTPUT: decode_62 
* OUTPUT: decode_63 
* OUTPUT: decode_64 
* OUTPUT: decode_65 
* OUTPUT: decode_66 
* OUTPUT: decode_67 
* OUTPUT: decode_68 
* OUTPUT: decode_69 
* OUTPUT: decode_70 
* OUTPUT: decode_71 
* OUTPUT: decode_72 
* OUTPUT: decode_73 
* OUTPUT: decode_74 
* OUTPUT: decode_75 
* OUTPUT: decode_76 
* OUTPUT: decode_77 
* OUTPUT: decode_78 
* OUTPUT: decode_79 
* OUTPUT: decode_80 
* OUTPUT: decode_81 
* OUTPUT: decode_82 
* OUTPUT: decode_83 
* OUTPUT: decode_84 
* OUTPUT: decode_85 
* OUTPUT: decode_86 
* OUTPUT: decode_87 
* OUTPUT: decode_88 
* OUTPUT: decode_89 
* OUTPUT: decode_90 
* OUTPUT: decode_91 
* OUTPUT: decode_92 
* OUTPUT: decode_93 
* OUTPUT: decode_94 
* OUTPUT: decode_95 
* OUTPUT: decode_96 
* OUTPUT: decode_97 
* OUTPUT: decode_98 
* OUTPUT: decode_99 
* OUTPUT: decode_100 
* OUTPUT: decode_101 
* OUTPUT: decode_102 
* OUTPUT: decode_103 
* OUTPUT: decode_104 
* OUTPUT: decode_105 
* OUTPUT: decode_106 
* OUTPUT: decode_107 
* OUTPUT: decode_108 
* OUTPUT: decode_109 
* OUTPUT: decode_110 
* OUTPUT: decode_111 
* OUTPUT: decode_112 
* OUTPUT: decode_113 
* OUTPUT: decode_114 
* OUTPUT: decode_115 
* OUTPUT: decode_116 
* OUTPUT: decode_117 
* OUTPUT: decode_118 
* OUTPUT: decode_119 
* OUTPUT: decode_120 
* OUTPUT: decode_121 
* OUTPUT: decode_122 
* OUTPUT: decode_123 
* OUTPUT: decode_124 
* OUTPUT: decode_125 
* OUTPUT: decode_126 
* OUTPUT: decode_127 
* OUTPUT: decode_128 
* POWER : vdd 
* GROUND: gnd 
Xpre_0 addr_0 addr_1 out_0 out_1 out_2 out_3 vdd gnd hierarchical_predecode2x4
Xpre3x8_0 addr_2 addr_3 addr_4 out_4 out_5 out_6 out_7 out_8 out_9 out_10 out_11 vdd gnd hierarchical_predecode3x8
Xpre3x8_1 addr_5 addr_6 addr_7 out_12 out_13 out_14 out_15 out_16 out_17 out_18 out_19 vdd gnd hierarchical_predecode3x8
XDEC_AND_0 out_0 out_4 out_12 decode_0 vdd gnd and3_dec
XDEC_AND_32 out_0 out_4 out_13 decode_32 vdd gnd and3_dec
XDEC_AND_64 out_0 out_4 out_14 decode_64 vdd gnd and3_dec
XDEC_AND_96 out_0 out_4 out_15 decode_96 vdd gnd and3_dec
XDEC_AND_128 out_0 out_4 out_16 decode_128 vdd gnd and3_dec
XDEC_AND_4 out_0 out_5 out_12 decode_4 vdd gnd and3_dec
XDEC_AND_36 out_0 out_5 out_13 decode_36 vdd gnd and3_dec
XDEC_AND_68 out_0 out_5 out_14 decode_68 vdd gnd and3_dec
XDEC_AND_100 out_0 out_5 out_15 decode_100 vdd gnd and3_dec
XDEC_AND_8 out_0 out_6 out_12 decode_8 vdd gnd and3_dec
XDEC_AND_40 out_0 out_6 out_13 decode_40 vdd gnd and3_dec
XDEC_AND_72 out_0 out_6 out_14 decode_72 vdd gnd and3_dec
XDEC_AND_104 out_0 out_6 out_15 decode_104 vdd gnd and3_dec
XDEC_AND_12 out_0 out_7 out_12 decode_12 vdd gnd and3_dec
XDEC_AND_44 out_0 out_7 out_13 decode_44 vdd gnd and3_dec
XDEC_AND_76 out_0 out_7 out_14 decode_76 vdd gnd and3_dec
XDEC_AND_108 out_0 out_7 out_15 decode_108 vdd gnd and3_dec
XDEC_AND_16 out_0 out_8 out_12 decode_16 vdd gnd and3_dec
XDEC_AND_48 out_0 out_8 out_13 decode_48 vdd gnd and3_dec
XDEC_AND_80 out_0 out_8 out_14 decode_80 vdd gnd and3_dec
XDEC_AND_112 out_0 out_8 out_15 decode_112 vdd gnd and3_dec
XDEC_AND_20 out_0 out_9 out_12 decode_20 vdd gnd and3_dec
XDEC_AND_52 out_0 out_9 out_13 decode_52 vdd gnd and3_dec
XDEC_AND_84 out_0 out_9 out_14 decode_84 vdd gnd and3_dec
XDEC_AND_116 out_0 out_9 out_15 decode_116 vdd gnd and3_dec
XDEC_AND_24 out_0 out_10 out_12 decode_24 vdd gnd and3_dec
XDEC_AND_56 out_0 out_10 out_13 decode_56 vdd gnd and3_dec
XDEC_AND_88 out_0 out_10 out_14 decode_88 vdd gnd and3_dec
XDEC_AND_120 out_0 out_10 out_15 decode_120 vdd gnd and3_dec
XDEC_AND_28 out_0 out_11 out_12 decode_28 vdd gnd and3_dec
XDEC_AND_60 out_0 out_11 out_13 decode_60 vdd gnd and3_dec
XDEC_AND_92 out_0 out_11 out_14 decode_92 vdd gnd and3_dec
XDEC_AND_124 out_0 out_11 out_15 decode_124 vdd gnd and3_dec
XDEC_AND_1 out_1 out_4 out_12 decode_1 vdd gnd and3_dec
XDEC_AND_33 out_1 out_4 out_13 decode_33 vdd gnd and3_dec
XDEC_AND_65 out_1 out_4 out_14 decode_65 vdd gnd and3_dec
XDEC_AND_97 out_1 out_4 out_15 decode_97 vdd gnd and3_dec
XDEC_AND_5 out_1 out_5 out_12 decode_5 vdd gnd and3_dec
XDEC_AND_37 out_1 out_5 out_13 decode_37 vdd gnd and3_dec
XDEC_AND_69 out_1 out_5 out_14 decode_69 vdd gnd and3_dec
XDEC_AND_101 out_1 out_5 out_15 decode_101 vdd gnd and3_dec
XDEC_AND_9 out_1 out_6 out_12 decode_9 vdd gnd and3_dec
XDEC_AND_41 out_1 out_6 out_13 decode_41 vdd gnd and3_dec
XDEC_AND_73 out_1 out_6 out_14 decode_73 vdd gnd and3_dec
XDEC_AND_105 out_1 out_6 out_15 decode_105 vdd gnd and3_dec
XDEC_AND_13 out_1 out_7 out_12 decode_13 vdd gnd and3_dec
XDEC_AND_45 out_1 out_7 out_13 decode_45 vdd gnd and3_dec
XDEC_AND_77 out_1 out_7 out_14 decode_77 vdd gnd and3_dec
XDEC_AND_109 out_1 out_7 out_15 decode_109 vdd gnd and3_dec
XDEC_AND_17 out_1 out_8 out_12 decode_17 vdd gnd and3_dec
XDEC_AND_49 out_1 out_8 out_13 decode_49 vdd gnd and3_dec
XDEC_AND_81 out_1 out_8 out_14 decode_81 vdd gnd and3_dec
XDEC_AND_113 out_1 out_8 out_15 decode_113 vdd gnd and3_dec
XDEC_AND_21 out_1 out_9 out_12 decode_21 vdd gnd and3_dec
XDEC_AND_53 out_1 out_9 out_13 decode_53 vdd gnd and3_dec
XDEC_AND_85 out_1 out_9 out_14 decode_85 vdd gnd and3_dec
XDEC_AND_117 out_1 out_9 out_15 decode_117 vdd gnd and3_dec
XDEC_AND_25 out_1 out_10 out_12 decode_25 vdd gnd and3_dec
XDEC_AND_57 out_1 out_10 out_13 decode_57 vdd gnd and3_dec
XDEC_AND_89 out_1 out_10 out_14 decode_89 vdd gnd and3_dec
XDEC_AND_121 out_1 out_10 out_15 decode_121 vdd gnd and3_dec
XDEC_AND_29 out_1 out_11 out_12 decode_29 vdd gnd and3_dec
XDEC_AND_61 out_1 out_11 out_13 decode_61 vdd gnd and3_dec
XDEC_AND_93 out_1 out_11 out_14 decode_93 vdd gnd and3_dec
XDEC_AND_125 out_1 out_11 out_15 decode_125 vdd gnd and3_dec
XDEC_AND_2 out_2 out_4 out_12 decode_2 vdd gnd and3_dec
XDEC_AND_34 out_2 out_4 out_13 decode_34 vdd gnd and3_dec
XDEC_AND_66 out_2 out_4 out_14 decode_66 vdd gnd and3_dec
XDEC_AND_98 out_2 out_4 out_15 decode_98 vdd gnd and3_dec
XDEC_AND_6 out_2 out_5 out_12 decode_6 vdd gnd and3_dec
XDEC_AND_38 out_2 out_5 out_13 decode_38 vdd gnd and3_dec
XDEC_AND_70 out_2 out_5 out_14 decode_70 vdd gnd and3_dec
XDEC_AND_102 out_2 out_5 out_15 decode_102 vdd gnd and3_dec
XDEC_AND_10 out_2 out_6 out_12 decode_10 vdd gnd and3_dec
XDEC_AND_42 out_2 out_6 out_13 decode_42 vdd gnd and3_dec
XDEC_AND_74 out_2 out_6 out_14 decode_74 vdd gnd and3_dec
XDEC_AND_106 out_2 out_6 out_15 decode_106 vdd gnd and3_dec
XDEC_AND_14 out_2 out_7 out_12 decode_14 vdd gnd and3_dec
XDEC_AND_46 out_2 out_7 out_13 decode_46 vdd gnd and3_dec
XDEC_AND_78 out_2 out_7 out_14 decode_78 vdd gnd and3_dec
XDEC_AND_110 out_2 out_7 out_15 decode_110 vdd gnd and3_dec
XDEC_AND_18 out_2 out_8 out_12 decode_18 vdd gnd and3_dec
XDEC_AND_50 out_2 out_8 out_13 decode_50 vdd gnd and3_dec
XDEC_AND_82 out_2 out_8 out_14 decode_82 vdd gnd and3_dec
XDEC_AND_114 out_2 out_8 out_15 decode_114 vdd gnd and3_dec
XDEC_AND_22 out_2 out_9 out_12 decode_22 vdd gnd and3_dec
XDEC_AND_54 out_2 out_9 out_13 decode_54 vdd gnd and3_dec
XDEC_AND_86 out_2 out_9 out_14 decode_86 vdd gnd and3_dec
XDEC_AND_118 out_2 out_9 out_15 decode_118 vdd gnd and3_dec
XDEC_AND_26 out_2 out_10 out_12 decode_26 vdd gnd and3_dec
XDEC_AND_58 out_2 out_10 out_13 decode_58 vdd gnd and3_dec
XDEC_AND_90 out_2 out_10 out_14 decode_90 vdd gnd and3_dec
XDEC_AND_122 out_2 out_10 out_15 decode_122 vdd gnd and3_dec
XDEC_AND_30 out_2 out_11 out_12 decode_30 vdd gnd and3_dec
XDEC_AND_62 out_2 out_11 out_13 decode_62 vdd gnd and3_dec
XDEC_AND_94 out_2 out_11 out_14 decode_94 vdd gnd and3_dec
XDEC_AND_126 out_2 out_11 out_15 decode_126 vdd gnd and3_dec
XDEC_AND_3 out_3 out_4 out_12 decode_3 vdd gnd and3_dec
XDEC_AND_35 out_3 out_4 out_13 decode_35 vdd gnd and3_dec
XDEC_AND_67 out_3 out_4 out_14 decode_67 vdd gnd and3_dec
XDEC_AND_99 out_3 out_4 out_15 decode_99 vdd gnd and3_dec
XDEC_AND_7 out_3 out_5 out_12 decode_7 vdd gnd and3_dec
XDEC_AND_39 out_3 out_5 out_13 decode_39 vdd gnd and3_dec
XDEC_AND_71 out_3 out_5 out_14 decode_71 vdd gnd and3_dec
XDEC_AND_103 out_3 out_5 out_15 decode_103 vdd gnd and3_dec
XDEC_AND_11 out_3 out_6 out_12 decode_11 vdd gnd and3_dec
XDEC_AND_43 out_3 out_6 out_13 decode_43 vdd gnd and3_dec
XDEC_AND_75 out_3 out_6 out_14 decode_75 vdd gnd and3_dec
XDEC_AND_107 out_3 out_6 out_15 decode_107 vdd gnd and3_dec
XDEC_AND_15 out_3 out_7 out_12 decode_15 vdd gnd and3_dec
XDEC_AND_47 out_3 out_7 out_13 decode_47 vdd gnd and3_dec
XDEC_AND_79 out_3 out_7 out_14 decode_79 vdd gnd and3_dec
XDEC_AND_111 out_3 out_7 out_15 decode_111 vdd gnd and3_dec
XDEC_AND_19 out_3 out_8 out_12 decode_19 vdd gnd and3_dec
XDEC_AND_51 out_3 out_8 out_13 decode_51 vdd gnd and3_dec
XDEC_AND_83 out_3 out_8 out_14 decode_83 vdd gnd and3_dec
XDEC_AND_115 out_3 out_8 out_15 decode_115 vdd gnd and3_dec
XDEC_AND_23 out_3 out_9 out_12 decode_23 vdd gnd and3_dec
XDEC_AND_55 out_3 out_9 out_13 decode_55 vdd gnd and3_dec
XDEC_AND_87 out_3 out_9 out_14 decode_87 vdd gnd and3_dec
XDEC_AND_119 out_3 out_9 out_15 decode_119 vdd gnd and3_dec
XDEC_AND_27 out_3 out_10 out_12 decode_27 vdd gnd and3_dec
XDEC_AND_59 out_3 out_10 out_13 decode_59 vdd gnd and3_dec
XDEC_AND_91 out_3 out_10 out_14 decode_91 vdd gnd and3_dec
XDEC_AND_123 out_3 out_10 out_15 decode_123 vdd gnd and3_dec
XDEC_AND_31 out_3 out_11 out_12 decode_31 vdd gnd and3_dec
XDEC_AND_63 out_3 out_11 out_13 decode_63 vdd gnd and3_dec
XDEC_AND_95 out_3 out_11 out_14 decode_95 vdd gnd and3_dec
XDEC_AND_127 out_3 out_11 out_15 decode_127 vdd gnd and3_dec
.ENDS hierarchical_decoder

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u

.SUBCKT pinv_dec_0 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
.ENDS pinv_dec_0

.SUBCKT wordline_driver A B Z vdd gnd
*.PININFO A:I B:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xwld_nand A B zb_int vdd gnd sky130_fd_bd_sram__openram_sp_nand2_dec
Xwl_driver zb_int Z vdd gnd pinv_dec_0
.ENDS wordline_driver

.SUBCKT wordline_driver_array in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12 in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23 in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34 in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45 in_46 in_47 in_48 in_49 in_50 in_51 in_52 in_53 in_54 in_55 in_56 in_57 in_58 in_59 in_60 in_61 in_62 in_63 in_64 in_65 in_66 in_67 in_68 in_69 in_70 in_71 in_72 in_73 in_74 in_75 in_76 in_77 in_78 in_79 in_80 in_81 in_82 in_83 in_84 in_85 in_86 in_87 in_88 in_89 in_90 in_91 in_92 in_93 in_94 in_95 in_96 in_97 in_98 in_99 in_100 in_101 in_102 in_103 in_104 in_105 in_106 in_107 in_108 in_109 in_110 in_111 in_112 in_113 in_114 in_115 in_116 in_117 in_118 in_119 in_120 in_121 in_122 in_123 in_124 in_125 in_126 in_127 in_128 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 en vdd gnd
*.PININFO in_0:I in_1:I in_2:I in_3:I in_4:I in_5:I in_6:I in_7:I in_8:I in_9:I in_10:I in_11:I in_12:I in_13:I in_14:I in_15:I in_16:I in_17:I in_18:I in_19:I in_20:I in_21:I in_22:I in_23:I in_24:I in_25:I in_26:I in_27:I in_28:I in_29:I in_30:I in_31:I in_32:I in_33:I in_34:I in_35:I in_36:I in_37:I in_38:I in_39:I in_40:I in_41:I in_42:I in_43:I in_44:I in_45:I in_46:I in_47:I in_48:I in_49:I in_50:I in_51:I in_52:I in_53:I in_54:I in_55:I in_56:I in_57:I in_58:I in_59:I in_60:I in_61:I in_62:I in_63:I in_64:I in_65:I in_66:I in_67:I in_68:I in_69:I in_70:I in_71:I in_72:I in_73:I in_74:I in_75:I in_76:I in_77:I in_78:I in_79:I in_80:I in_81:I in_82:I in_83:I in_84:I in_85:I in_86:I in_87:I in_88:I in_89:I in_90:I in_91:I in_92:I in_93:I in_94:I in_95:I in_96:I in_97:I in_98:I in_99:I in_100:I in_101:I in_102:I in_103:I in_104:I in_105:I in_106:I in_107:I in_108:I in_109:I in_110:I in_111:I in_112:I in_113:I in_114:I in_115:I in_116:I in_117:I in_118:I in_119:I in_120:I in_121:I in_122:I in_123:I in_124:I in_125:I in_126:I in_127:I in_128:I wl_0:O wl_1:O wl_2:O wl_3:O wl_4:O wl_5:O wl_6:O wl_7:O wl_8:O wl_9:O wl_10:O wl_11:O wl_12:O wl_13:O wl_14:O wl_15:O wl_16:O wl_17:O wl_18:O wl_19:O wl_20:O wl_21:O wl_22:O wl_23:O wl_24:O wl_25:O wl_26:O wl_27:O wl_28:O wl_29:O wl_30:O wl_31:O wl_32:O wl_33:O wl_34:O wl_35:O wl_36:O wl_37:O wl_38:O wl_39:O wl_40:O wl_41:O wl_42:O wl_43:O wl_44:O wl_45:O wl_46:O wl_47:O wl_48:O wl_49:O wl_50:O wl_51:O wl_52:O wl_53:O wl_54:O wl_55:O wl_56:O wl_57:O wl_58:O wl_59:O wl_60:O wl_61:O wl_62:O wl_63:O wl_64:O wl_65:O wl_66:O wl_67:O wl_68:O wl_69:O wl_70:O wl_71:O wl_72:O wl_73:O wl_74:O wl_75:O wl_76:O wl_77:O wl_78:O wl_79:O wl_80:O wl_81:O wl_82:O wl_83:O wl_84:O wl_85:O wl_86:O wl_87:O wl_88:O wl_89:O wl_90:O wl_91:O wl_92:O wl_93:O wl_94:O wl_95:O wl_96:O wl_97:O wl_98:O wl_99:O wl_100:O wl_101:O wl_102:O wl_103:O wl_104:O wl_105:O wl_106:O wl_107:O wl_108:O wl_109:O wl_110:O wl_111:O wl_112:O wl_113:O wl_114:O wl_115:O wl_116:O wl_117:O wl_118:O wl_119:O wl_120:O wl_121:O wl_122:O wl_123:O wl_124:O wl_125:O wl_126:O wl_127:O wl_128:O en:I vdd:B gnd:B
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* INPUT : in_32 
* INPUT : in_33 
* INPUT : in_34 
* INPUT : in_35 
* INPUT : in_36 
* INPUT : in_37 
* INPUT : in_38 
* INPUT : in_39 
* INPUT : in_40 
* INPUT : in_41 
* INPUT : in_42 
* INPUT : in_43 
* INPUT : in_44 
* INPUT : in_45 
* INPUT : in_46 
* INPUT : in_47 
* INPUT : in_48 
* INPUT : in_49 
* INPUT : in_50 
* INPUT : in_51 
* INPUT : in_52 
* INPUT : in_53 
* INPUT : in_54 
* INPUT : in_55 
* INPUT : in_56 
* INPUT : in_57 
* INPUT : in_58 
* INPUT : in_59 
* INPUT : in_60 
* INPUT : in_61 
* INPUT : in_62 
* INPUT : in_63 
* INPUT : in_64 
* INPUT : in_65 
* INPUT : in_66 
* INPUT : in_67 
* INPUT : in_68 
* INPUT : in_69 
* INPUT : in_70 
* INPUT : in_71 
* INPUT : in_72 
* INPUT : in_73 
* INPUT : in_74 
* INPUT : in_75 
* INPUT : in_76 
* INPUT : in_77 
* INPUT : in_78 
* INPUT : in_79 
* INPUT : in_80 
* INPUT : in_81 
* INPUT : in_82 
* INPUT : in_83 
* INPUT : in_84 
* INPUT : in_85 
* INPUT : in_86 
* INPUT : in_87 
* INPUT : in_88 
* INPUT : in_89 
* INPUT : in_90 
* INPUT : in_91 
* INPUT : in_92 
* INPUT : in_93 
* INPUT : in_94 
* INPUT : in_95 
* INPUT : in_96 
* INPUT : in_97 
* INPUT : in_98 
* INPUT : in_99 
* INPUT : in_100 
* INPUT : in_101 
* INPUT : in_102 
* INPUT : in_103 
* INPUT : in_104 
* INPUT : in_105 
* INPUT : in_106 
* INPUT : in_107 
* INPUT : in_108 
* INPUT : in_109 
* INPUT : in_110 
* INPUT : in_111 
* INPUT : in_112 
* INPUT : in_113 
* INPUT : in_114 
* INPUT : in_115 
* INPUT : in_116 
* INPUT : in_117 
* INPUT : in_118 
* INPUT : in_119 
* INPUT : in_120 
* INPUT : in_121 
* INPUT : in_122 
* INPUT : in_123 
* INPUT : in_124 
* INPUT : in_125 
* INPUT : in_126 
* INPUT : in_127 
* INPUT : in_128 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* OUTPUT: wl_89 
* OUTPUT: wl_90 
* OUTPUT: wl_91 
* OUTPUT: wl_92 
* OUTPUT: wl_93 
* OUTPUT: wl_94 
* OUTPUT: wl_95 
* OUTPUT: wl_96 
* OUTPUT: wl_97 
* OUTPUT: wl_98 
* OUTPUT: wl_99 
* OUTPUT: wl_100 
* OUTPUT: wl_101 
* OUTPUT: wl_102 
* OUTPUT: wl_103 
* OUTPUT: wl_104 
* OUTPUT: wl_105 
* OUTPUT: wl_106 
* OUTPUT: wl_107 
* OUTPUT: wl_108 
* OUTPUT: wl_109 
* OUTPUT: wl_110 
* OUTPUT: wl_111 
* OUTPUT: wl_112 
* OUTPUT: wl_113 
* OUTPUT: wl_114 
* OUTPUT: wl_115 
* OUTPUT: wl_116 
* OUTPUT: wl_117 
* OUTPUT: wl_118 
* OUTPUT: wl_119 
* OUTPUT: wl_120 
* OUTPUT: wl_121 
* OUTPUT: wl_122 
* OUTPUT: wl_123 
* OUTPUT: wl_124 
* OUTPUT: wl_125 
* OUTPUT: wl_126 
* OUTPUT: wl_127 
* OUTPUT: wl_128 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* rows: 129 cols: 129
Xwl_driver_and0 in_0 en wl_0 vdd gnd wordline_driver
Xwl_driver_and1 in_1 en wl_1 vdd gnd wordline_driver
Xwl_driver_and2 in_2 en wl_2 vdd gnd wordline_driver
Xwl_driver_and3 in_3 en wl_3 vdd gnd wordline_driver
Xwl_driver_and4 in_4 en wl_4 vdd gnd wordline_driver
Xwl_driver_and5 in_5 en wl_5 vdd gnd wordline_driver
Xwl_driver_and6 in_6 en wl_6 vdd gnd wordline_driver
Xwl_driver_and7 in_7 en wl_7 vdd gnd wordline_driver
Xwl_driver_and8 in_8 en wl_8 vdd gnd wordline_driver
Xwl_driver_and9 in_9 en wl_9 vdd gnd wordline_driver
Xwl_driver_and10 in_10 en wl_10 vdd gnd wordline_driver
Xwl_driver_and11 in_11 en wl_11 vdd gnd wordline_driver
Xwl_driver_and12 in_12 en wl_12 vdd gnd wordline_driver
Xwl_driver_and13 in_13 en wl_13 vdd gnd wordline_driver
Xwl_driver_and14 in_14 en wl_14 vdd gnd wordline_driver
Xwl_driver_and15 in_15 en wl_15 vdd gnd wordline_driver
Xwl_driver_and16 in_16 en wl_16 vdd gnd wordline_driver
Xwl_driver_and17 in_17 en wl_17 vdd gnd wordline_driver
Xwl_driver_and18 in_18 en wl_18 vdd gnd wordline_driver
Xwl_driver_and19 in_19 en wl_19 vdd gnd wordline_driver
Xwl_driver_and20 in_20 en wl_20 vdd gnd wordline_driver
Xwl_driver_and21 in_21 en wl_21 vdd gnd wordline_driver
Xwl_driver_and22 in_22 en wl_22 vdd gnd wordline_driver
Xwl_driver_and23 in_23 en wl_23 vdd gnd wordline_driver
Xwl_driver_and24 in_24 en wl_24 vdd gnd wordline_driver
Xwl_driver_and25 in_25 en wl_25 vdd gnd wordline_driver
Xwl_driver_and26 in_26 en wl_26 vdd gnd wordline_driver
Xwl_driver_and27 in_27 en wl_27 vdd gnd wordline_driver
Xwl_driver_and28 in_28 en wl_28 vdd gnd wordline_driver
Xwl_driver_and29 in_29 en wl_29 vdd gnd wordline_driver
Xwl_driver_and30 in_30 en wl_30 vdd gnd wordline_driver
Xwl_driver_and31 in_31 en wl_31 vdd gnd wordline_driver
Xwl_driver_and32 in_32 en wl_32 vdd gnd wordline_driver
Xwl_driver_and33 in_33 en wl_33 vdd gnd wordline_driver
Xwl_driver_and34 in_34 en wl_34 vdd gnd wordline_driver
Xwl_driver_and35 in_35 en wl_35 vdd gnd wordline_driver
Xwl_driver_and36 in_36 en wl_36 vdd gnd wordline_driver
Xwl_driver_and37 in_37 en wl_37 vdd gnd wordline_driver
Xwl_driver_and38 in_38 en wl_38 vdd gnd wordline_driver
Xwl_driver_and39 in_39 en wl_39 vdd gnd wordline_driver
Xwl_driver_and40 in_40 en wl_40 vdd gnd wordline_driver
Xwl_driver_and41 in_41 en wl_41 vdd gnd wordline_driver
Xwl_driver_and42 in_42 en wl_42 vdd gnd wordline_driver
Xwl_driver_and43 in_43 en wl_43 vdd gnd wordline_driver
Xwl_driver_and44 in_44 en wl_44 vdd gnd wordline_driver
Xwl_driver_and45 in_45 en wl_45 vdd gnd wordline_driver
Xwl_driver_and46 in_46 en wl_46 vdd gnd wordline_driver
Xwl_driver_and47 in_47 en wl_47 vdd gnd wordline_driver
Xwl_driver_and48 in_48 en wl_48 vdd gnd wordline_driver
Xwl_driver_and49 in_49 en wl_49 vdd gnd wordline_driver
Xwl_driver_and50 in_50 en wl_50 vdd gnd wordline_driver
Xwl_driver_and51 in_51 en wl_51 vdd gnd wordline_driver
Xwl_driver_and52 in_52 en wl_52 vdd gnd wordline_driver
Xwl_driver_and53 in_53 en wl_53 vdd gnd wordline_driver
Xwl_driver_and54 in_54 en wl_54 vdd gnd wordline_driver
Xwl_driver_and55 in_55 en wl_55 vdd gnd wordline_driver
Xwl_driver_and56 in_56 en wl_56 vdd gnd wordline_driver
Xwl_driver_and57 in_57 en wl_57 vdd gnd wordline_driver
Xwl_driver_and58 in_58 en wl_58 vdd gnd wordline_driver
Xwl_driver_and59 in_59 en wl_59 vdd gnd wordline_driver
Xwl_driver_and60 in_60 en wl_60 vdd gnd wordline_driver
Xwl_driver_and61 in_61 en wl_61 vdd gnd wordline_driver
Xwl_driver_and62 in_62 en wl_62 vdd gnd wordline_driver
Xwl_driver_and63 in_63 en wl_63 vdd gnd wordline_driver
Xwl_driver_and64 in_64 en wl_64 vdd gnd wordline_driver
Xwl_driver_and65 in_65 en wl_65 vdd gnd wordline_driver
Xwl_driver_and66 in_66 en wl_66 vdd gnd wordline_driver
Xwl_driver_and67 in_67 en wl_67 vdd gnd wordline_driver
Xwl_driver_and68 in_68 en wl_68 vdd gnd wordline_driver
Xwl_driver_and69 in_69 en wl_69 vdd gnd wordline_driver
Xwl_driver_and70 in_70 en wl_70 vdd gnd wordline_driver
Xwl_driver_and71 in_71 en wl_71 vdd gnd wordline_driver
Xwl_driver_and72 in_72 en wl_72 vdd gnd wordline_driver
Xwl_driver_and73 in_73 en wl_73 vdd gnd wordline_driver
Xwl_driver_and74 in_74 en wl_74 vdd gnd wordline_driver
Xwl_driver_and75 in_75 en wl_75 vdd gnd wordline_driver
Xwl_driver_and76 in_76 en wl_76 vdd gnd wordline_driver
Xwl_driver_and77 in_77 en wl_77 vdd gnd wordline_driver
Xwl_driver_and78 in_78 en wl_78 vdd gnd wordline_driver
Xwl_driver_and79 in_79 en wl_79 vdd gnd wordline_driver
Xwl_driver_and80 in_80 en wl_80 vdd gnd wordline_driver
Xwl_driver_and81 in_81 en wl_81 vdd gnd wordline_driver
Xwl_driver_and82 in_82 en wl_82 vdd gnd wordline_driver
Xwl_driver_and83 in_83 en wl_83 vdd gnd wordline_driver
Xwl_driver_and84 in_84 en wl_84 vdd gnd wordline_driver
Xwl_driver_and85 in_85 en wl_85 vdd gnd wordline_driver
Xwl_driver_and86 in_86 en wl_86 vdd gnd wordline_driver
Xwl_driver_and87 in_87 en wl_87 vdd gnd wordline_driver
Xwl_driver_and88 in_88 en wl_88 vdd gnd wordline_driver
Xwl_driver_and89 in_89 en wl_89 vdd gnd wordline_driver
Xwl_driver_and90 in_90 en wl_90 vdd gnd wordline_driver
Xwl_driver_and91 in_91 en wl_91 vdd gnd wordline_driver
Xwl_driver_and92 in_92 en wl_92 vdd gnd wordline_driver
Xwl_driver_and93 in_93 en wl_93 vdd gnd wordline_driver
Xwl_driver_and94 in_94 en wl_94 vdd gnd wordline_driver
Xwl_driver_and95 in_95 en wl_95 vdd gnd wordline_driver
Xwl_driver_and96 in_96 en wl_96 vdd gnd wordline_driver
Xwl_driver_and97 in_97 en wl_97 vdd gnd wordline_driver
Xwl_driver_and98 in_98 en wl_98 vdd gnd wordline_driver
Xwl_driver_and99 in_99 en wl_99 vdd gnd wordline_driver
Xwl_driver_and100 in_100 en wl_100 vdd gnd wordline_driver
Xwl_driver_and101 in_101 en wl_101 vdd gnd wordline_driver
Xwl_driver_and102 in_102 en wl_102 vdd gnd wordline_driver
Xwl_driver_and103 in_103 en wl_103 vdd gnd wordline_driver
Xwl_driver_and104 in_104 en wl_104 vdd gnd wordline_driver
Xwl_driver_and105 in_105 en wl_105 vdd gnd wordline_driver
Xwl_driver_and106 in_106 en wl_106 vdd gnd wordline_driver
Xwl_driver_and107 in_107 en wl_107 vdd gnd wordline_driver
Xwl_driver_and108 in_108 en wl_108 vdd gnd wordline_driver
Xwl_driver_and109 in_109 en wl_109 vdd gnd wordline_driver
Xwl_driver_and110 in_110 en wl_110 vdd gnd wordline_driver
Xwl_driver_and111 in_111 en wl_111 vdd gnd wordline_driver
Xwl_driver_and112 in_112 en wl_112 vdd gnd wordline_driver
Xwl_driver_and113 in_113 en wl_113 vdd gnd wordline_driver
Xwl_driver_and114 in_114 en wl_114 vdd gnd wordline_driver
Xwl_driver_and115 in_115 en wl_115 vdd gnd wordline_driver
Xwl_driver_and116 in_116 en wl_116 vdd gnd wordline_driver
Xwl_driver_and117 in_117 en wl_117 vdd gnd wordline_driver
Xwl_driver_and118 in_118 en wl_118 vdd gnd wordline_driver
Xwl_driver_and119 in_119 en wl_119 vdd gnd wordline_driver
Xwl_driver_and120 in_120 en wl_120 vdd gnd wordline_driver
Xwl_driver_and121 in_121 en wl_121 vdd gnd wordline_driver
Xwl_driver_and122 in_122 en wl_122 vdd gnd wordline_driver
Xwl_driver_and123 in_123 en wl_123 vdd gnd wordline_driver
Xwl_driver_and124 in_124 en wl_124 vdd gnd wordline_driver
Xwl_driver_and125 in_125 en wl_125 vdd gnd wordline_driver
Xwl_driver_and126 in_126 en wl_126 vdd gnd wordline_driver
Xwl_driver_and127 in_127 en wl_127 vdd gnd wordline_driver
Xwl_driver_and128 in_128 en wl_128 vdd gnd wordline_driver
.ENDS wordline_driver_array

.SUBCKT and2_dec_0 A B Z vdd gnd
*.PININFO A:I B:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 32
Xpand2_dec_nand A B zb_int vdd gnd sky130_fd_bd_sram__openram_sp_nand2_dec
Xpand2_dec_inv zb_int Z vdd gnd pinv_dec_0
.ENDS and2_dec_0

.SUBCKT port_address addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 addr_7 wl_en wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 rbl_wl vdd gnd
*.PININFO addr_0:I addr_1:I addr_2:I addr_3:I addr_4:I addr_5:I addr_6:I addr_7:I wl_en:I wl_0:O wl_1:O wl_2:O wl_3:O wl_4:O wl_5:O wl_6:O wl_7:O wl_8:O wl_9:O wl_10:O wl_11:O wl_12:O wl_13:O wl_14:O wl_15:O wl_16:O wl_17:O wl_18:O wl_19:O wl_20:O wl_21:O wl_22:O wl_23:O wl_24:O wl_25:O wl_26:O wl_27:O wl_28:O wl_29:O wl_30:O wl_31:O wl_32:O wl_33:O wl_34:O wl_35:O wl_36:O wl_37:O wl_38:O wl_39:O wl_40:O wl_41:O wl_42:O wl_43:O wl_44:O wl_45:O wl_46:O wl_47:O wl_48:O wl_49:O wl_50:O wl_51:O wl_52:O wl_53:O wl_54:O wl_55:O wl_56:O wl_57:O wl_58:O wl_59:O wl_60:O wl_61:O wl_62:O wl_63:O wl_64:O wl_65:O wl_66:O wl_67:O wl_68:O wl_69:O wl_70:O wl_71:O wl_72:O wl_73:O wl_74:O wl_75:O wl_76:O wl_77:O wl_78:O wl_79:O wl_80:O wl_81:O wl_82:O wl_83:O wl_84:O wl_85:O wl_86:O wl_87:O wl_88:O wl_89:O wl_90:O wl_91:O wl_92:O wl_93:O wl_94:O wl_95:O wl_96:O wl_97:O wl_98:O wl_99:O wl_100:O wl_101:O wl_102:O wl_103:O wl_104:O wl_105:O wl_106:O wl_107:O wl_108:O wl_109:O wl_110:O wl_111:O wl_112:O wl_113:O wl_114:O wl_115:O wl_116:O wl_117:O wl_118:O wl_119:O wl_120:O wl_121:O wl_122:O wl_123:O wl_124:O wl_125:O wl_126:O wl_127:O wl_128:O rbl_wl:O vdd:B gnd:B
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* INPUT : addr_7 
* INPUT : wl_en 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* OUTPUT: wl_89 
* OUTPUT: wl_90 
* OUTPUT: wl_91 
* OUTPUT: wl_92 
* OUTPUT: wl_93 
* OUTPUT: wl_94 
* OUTPUT: wl_95 
* OUTPUT: wl_96 
* OUTPUT: wl_97 
* OUTPUT: wl_98 
* OUTPUT: wl_99 
* OUTPUT: wl_100 
* OUTPUT: wl_101 
* OUTPUT: wl_102 
* OUTPUT: wl_103 
* OUTPUT: wl_104 
* OUTPUT: wl_105 
* OUTPUT: wl_106 
* OUTPUT: wl_107 
* OUTPUT: wl_108 
* OUTPUT: wl_109 
* OUTPUT: wl_110 
* OUTPUT: wl_111 
* OUTPUT: wl_112 
* OUTPUT: wl_113 
* OUTPUT: wl_114 
* OUTPUT: wl_115 
* OUTPUT: wl_116 
* OUTPUT: wl_117 
* OUTPUT: wl_118 
* OUTPUT: wl_119 
* OUTPUT: wl_120 
* OUTPUT: wl_121 
* OUTPUT: wl_122 
* OUTPUT: wl_123 
* OUTPUT: wl_124 
* OUTPUT: wl_125 
* OUTPUT: wl_126 
* OUTPUT: wl_127 
* OUTPUT: wl_128 
* OUTPUT: rbl_wl 
* POWER : vdd 
* GROUND: gnd 
Xrow_decoder addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 addr_7 dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62 dec_out_63 dec_out_64 dec_out_65 dec_out_66 dec_out_67 dec_out_68 dec_out_69 dec_out_70 dec_out_71 dec_out_72 dec_out_73 dec_out_74 dec_out_75 dec_out_76 dec_out_77 dec_out_78 dec_out_79 dec_out_80 dec_out_81 dec_out_82 dec_out_83 dec_out_84 dec_out_85 dec_out_86 dec_out_87 dec_out_88 dec_out_89 dec_out_90 dec_out_91 dec_out_92 dec_out_93 dec_out_94 dec_out_95 dec_out_96 dec_out_97 dec_out_98 dec_out_99 dec_out_100 dec_out_101 dec_out_102 dec_out_103 dec_out_104 dec_out_105 dec_out_106 dec_out_107 dec_out_108 dec_out_109 dec_out_110 dec_out_111 dec_out_112 dec_out_113 dec_out_114 dec_out_115 dec_out_116 dec_out_117 dec_out_118 dec_out_119 dec_out_120 dec_out_121 dec_out_122 dec_out_123 dec_out_124 dec_out_125 dec_out_126 dec_out_127 dec_out_128 vdd gnd hierarchical_decoder
Xwordline_driver dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62 dec_out_63 dec_out_64 dec_out_65 dec_out_66 dec_out_67 dec_out_68 dec_out_69 dec_out_70 dec_out_71 dec_out_72 dec_out_73 dec_out_74 dec_out_75 dec_out_76 dec_out_77 dec_out_78 dec_out_79 dec_out_80 dec_out_81 dec_out_82 dec_out_83 dec_out_84 dec_out_85 dec_out_86 dec_out_87 dec_out_88 dec_out_89 dec_out_90 dec_out_91 dec_out_92 dec_out_93 dec_out_94 dec_out_95 dec_out_96 dec_out_97 dec_out_98 dec_out_99 dec_out_100 dec_out_101 dec_out_102 dec_out_103 dec_out_104 dec_out_105 dec_out_106 dec_out_107 dec_out_108 dec_out_109 dec_out_110 dec_out_111 dec_out_112 dec_out_113 dec_out_114 dec_out_115 dec_out_116 dec_out_117 dec_out_118 dec_out_119 dec_out_120 dec_out_121 dec_out_122 dec_out_123 dec_out_124 dec_out_125 dec_out_126 dec_out_127 dec_out_128 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_en vdd gnd wordline_driver_array
Xrbl_driver wl_en vdd rbl_wl vdd gnd and2_dec_0
.ENDS port_address

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u

.SUBCKT precharge_0 bl br en_bar vdd
*.PININFO bl:O br:O en_bar:I vdd:B
* OUTPUT: bl 
* OUTPUT: br 
* INPUT : en_bar 
* POWER : vdd 
Xlower_pmos bl en_bar br vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
Xupper_pmos1 bl en_bar vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
Xupper_pmos2 br en_bar vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
.ENDS precharge_0

.SUBCKT precharge_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 en_bar vdd
*.PININFO bl_0:O br_0:O bl_1:O br_1:O bl_2:O br_2:O bl_3:O br_3:O bl_4:O br_4:O bl_5:O br_5:O bl_6:O br_6:O bl_7:O br_7:O bl_8:O br_8:O bl_9:O br_9:O bl_10:O br_10:O bl_11:O br_11:O bl_12:O br_12:O bl_13:O br_13:O bl_14:O br_14:O bl_15:O br_15:O bl_16:O br_16:O bl_17:O br_17:O bl_18:O br_18:O bl_19:O br_19:O bl_20:O br_20:O bl_21:O br_21:O bl_22:O br_22:O bl_23:O br_23:O bl_24:O br_24:O bl_25:O br_25:O bl_26:O br_26:O bl_27:O br_27:O bl_28:O br_28:O bl_29:O br_29:O bl_30:O br_30:O bl_31:O br_31:O bl_32:O br_32:O bl_33:O br_33:O bl_34:O br_34:O bl_35:O br_35:O bl_36:O br_36:O bl_37:O br_37:O bl_38:O br_38:O bl_39:O br_39:O bl_40:O br_40:O bl_41:O br_41:O bl_42:O br_42:O bl_43:O br_43:O bl_44:O br_44:O bl_45:O br_45:O bl_46:O br_46:O bl_47:O br_47:O bl_48:O br_48:O bl_49:O br_49:O bl_50:O br_50:O bl_51:O br_51:O bl_52:O br_52:O bl_53:O br_53:O bl_54:O br_54:O bl_55:O br_55:O bl_56:O br_56:O bl_57:O br_57:O bl_58:O br_58:O bl_59:O br_59:O bl_60:O br_60:O bl_61:O br_61:O bl_62:O br_62:O bl_63:O br_63:O bl_64:O br_64:O bl_65:O br_65:O bl_66:O br_66:O bl_67:O br_67:O bl_68:O br_68:O bl_69:O br_69:O bl_70:O br_70:O bl_71:O br_71:O bl_72:O br_72:O bl_73:O br_73:O bl_74:O br_74:O bl_75:O br_75:O bl_76:O br_76:O bl_77:O br_77:O bl_78:O br_78:O bl_79:O br_79:O bl_80:O br_80:O bl_81:O br_81:O bl_82:O br_82:O bl_83:O br_83:O bl_84:O br_84:O bl_85:O br_85:O bl_86:O br_86:O bl_87:O br_87:O bl_88:O br_88:O bl_89:O br_89:O bl_90:O br_90:O bl_91:O br_91:O bl_92:O br_92:O bl_93:O br_93:O bl_94:O br_94:O bl_95:O br_95:O bl_96:O br_96:O bl_97:O br_97:O bl_98:O br_98:O bl_99:O br_99:O bl_100:O br_100:O bl_101:O br_101:O bl_102:O br_102:O bl_103:O br_103:O bl_104:O br_104:O bl_105:O br_105:O bl_106:O br_106:O bl_107:O br_107:O bl_108:O br_108:O bl_109:O br_109:O bl_110:O br_110:O bl_111:O br_111:O bl_112:O br_112:O bl_113:O br_113:O bl_114:O br_114:O bl_115:O br_115:O bl_116:O br_116:O bl_117:O br_117:O bl_118:O br_118:O bl_119:O br_119:O bl_120:O br_120:O bl_121:O br_121:O bl_122:O br_122:O bl_123:O br_123:O bl_124:O br_124:O bl_125:O br_125:O bl_126:O br_126:O bl_127:O br_127:O bl_128:O br_128:O bl_129:O br_129:O en_bar:I vdd:B
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* OUTPUT: bl_65 
* OUTPUT: br_65 
* OUTPUT: bl_66 
* OUTPUT: br_66 
* OUTPUT: bl_67 
* OUTPUT: br_67 
* OUTPUT: bl_68 
* OUTPUT: br_68 
* OUTPUT: bl_69 
* OUTPUT: br_69 
* OUTPUT: bl_70 
* OUTPUT: br_70 
* OUTPUT: bl_71 
* OUTPUT: br_71 
* OUTPUT: bl_72 
* OUTPUT: br_72 
* OUTPUT: bl_73 
* OUTPUT: br_73 
* OUTPUT: bl_74 
* OUTPUT: br_74 
* OUTPUT: bl_75 
* OUTPUT: br_75 
* OUTPUT: bl_76 
* OUTPUT: br_76 
* OUTPUT: bl_77 
* OUTPUT: br_77 
* OUTPUT: bl_78 
* OUTPUT: br_78 
* OUTPUT: bl_79 
* OUTPUT: br_79 
* OUTPUT: bl_80 
* OUTPUT: br_80 
* OUTPUT: bl_81 
* OUTPUT: br_81 
* OUTPUT: bl_82 
* OUTPUT: br_82 
* OUTPUT: bl_83 
* OUTPUT: br_83 
* OUTPUT: bl_84 
* OUTPUT: br_84 
* OUTPUT: bl_85 
* OUTPUT: br_85 
* OUTPUT: bl_86 
* OUTPUT: br_86 
* OUTPUT: bl_87 
* OUTPUT: br_87 
* OUTPUT: bl_88 
* OUTPUT: br_88 
* OUTPUT: bl_89 
* OUTPUT: br_89 
* OUTPUT: bl_90 
* OUTPUT: br_90 
* OUTPUT: bl_91 
* OUTPUT: br_91 
* OUTPUT: bl_92 
* OUTPUT: br_92 
* OUTPUT: bl_93 
* OUTPUT: br_93 
* OUTPUT: bl_94 
* OUTPUT: br_94 
* OUTPUT: bl_95 
* OUTPUT: br_95 
* OUTPUT: bl_96 
* OUTPUT: br_96 
* OUTPUT: bl_97 
* OUTPUT: br_97 
* OUTPUT: bl_98 
* OUTPUT: br_98 
* OUTPUT: bl_99 
* OUTPUT: br_99 
* OUTPUT: bl_100 
* OUTPUT: br_100 
* OUTPUT: bl_101 
* OUTPUT: br_101 
* OUTPUT: bl_102 
* OUTPUT: br_102 
* OUTPUT: bl_103 
* OUTPUT: br_103 
* OUTPUT: bl_104 
* OUTPUT: br_104 
* OUTPUT: bl_105 
* OUTPUT: br_105 
* OUTPUT: bl_106 
* OUTPUT: br_106 
* OUTPUT: bl_107 
* OUTPUT: br_107 
* OUTPUT: bl_108 
* OUTPUT: br_108 
* OUTPUT: bl_109 
* OUTPUT: br_109 
* OUTPUT: bl_110 
* OUTPUT: br_110 
* OUTPUT: bl_111 
* OUTPUT: br_111 
* OUTPUT: bl_112 
* OUTPUT: br_112 
* OUTPUT: bl_113 
* OUTPUT: br_113 
* OUTPUT: bl_114 
* OUTPUT: br_114 
* OUTPUT: bl_115 
* OUTPUT: br_115 
* OUTPUT: bl_116 
* OUTPUT: br_116 
* OUTPUT: bl_117 
* OUTPUT: br_117 
* OUTPUT: bl_118 
* OUTPUT: br_118 
* OUTPUT: bl_119 
* OUTPUT: br_119 
* OUTPUT: bl_120 
* OUTPUT: br_120 
* OUTPUT: bl_121 
* OUTPUT: br_121 
* OUTPUT: bl_122 
* OUTPUT: br_122 
* OUTPUT: bl_123 
* OUTPUT: br_123 
* OUTPUT: bl_124 
* OUTPUT: br_124 
* OUTPUT: bl_125 
* OUTPUT: br_125 
* OUTPUT: bl_126 
* OUTPUT: br_126 
* OUTPUT: bl_127 
* OUTPUT: br_127 
* OUTPUT: bl_128 
* OUTPUT: br_128 
* OUTPUT: bl_129 
* OUTPUT: br_129 
* INPUT : en_bar 
* POWER : vdd 
* cols: 130 size: 1 bl: bl br: br
Xpre_column_0 bl_0 br_0 en_bar vdd precharge_0
Xpre_column_1 bl_1 br_1 en_bar vdd precharge_0
Xpre_column_2 bl_2 br_2 en_bar vdd precharge_0
Xpre_column_3 bl_3 br_3 en_bar vdd precharge_0
Xpre_column_4 bl_4 br_4 en_bar vdd precharge_0
Xpre_column_5 bl_5 br_5 en_bar vdd precharge_0
Xpre_column_6 bl_6 br_6 en_bar vdd precharge_0
Xpre_column_7 bl_7 br_7 en_bar vdd precharge_0
Xpre_column_8 bl_8 br_8 en_bar vdd precharge_0
Xpre_column_9 bl_9 br_9 en_bar vdd precharge_0
Xpre_column_10 bl_10 br_10 en_bar vdd precharge_0
Xpre_column_11 bl_11 br_11 en_bar vdd precharge_0
Xpre_column_12 bl_12 br_12 en_bar vdd precharge_0
Xpre_column_13 bl_13 br_13 en_bar vdd precharge_0
Xpre_column_14 bl_14 br_14 en_bar vdd precharge_0
Xpre_column_15 bl_15 br_15 en_bar vdd precharge_0
Xpre_column_16 bl_16 br_16 en_bar vdd precharge_0
Xpre_column_17 bl_17 br_17 en_bar vdd precharge_0
Xpre_column_18 bl_18 br_18 en_bar vdd precharge_0
Xpre_column_19 bl_19 br_19 en_bar vdd precharge_0
Xpre_column_20 bl_20 br_20 en_bar vdd precharge_0
Xpre_column_21 bl_21 br_21 en_bar vdd precharge_0
Xpre_column_22 bl_22 br_22 en_bar vdd precharge_0
Xpre_column_23 bl_23 br_23 en_bar vdd precharge_0
Xpre_column_24 bl_24 br_24 en_bar vdd precharge_0
Xpre_column_25 bl_25 br_25 en_bar vdd precharge_0
Xpre_column_26 bl_26 br_26 en_bar vdd precharge_0
Xpre_column_27 bl_27 br_27 en_bar vdd precharge_0
Xpre_column_28 bl_28 br_28 en_bar vdd precharge_0
Xpre_column_29 bl_29 br_29 en_bar vdd precharge_0
Xpre_column_30 bl_30 br_30 en_bar vdd precharge_0
Xpre_column_31 bl_31 br_31 en_bar vdd precharge_0
Xpre_column_32 bl_32 br_32 en_bar vdd precharge_0
Xpre_column_33 bl_33 br_33 en_bar vdd precharge_0
Xpre_column_34 bl_34 br_34 en_bar vdd precharge_0
Xpre_column_35 bl_35 br_35 en_bar vdd precharge_0
Xpre_column_36 bl_36 br_36 en_bar vdd precharge_0
Xpre_column_37 bl_37 br_37 en_bar vdd precharge_0
Xpre_column_38 bl_38 br_38 en_bar vdd precharge_0
Xpre_column_39 bl_39 br_39 en_bar vdd precharge_0
Xpre_column_40 bl_40 br_40 en_bar vdd precharge_0
Xpre_column_41 bl_41 br_41 en_bar vdd precharge_0
Xpre_column_42 bl_42 br_42 en_bar vdd precharge_0
Xpre_column_43 bl_43 br_43 en_bar vdd precharge_0
Xpre_column_44 bl_44 br_44 en_bar vdd precharge_0
Xpre_column_45 bl_45 br_45 en_bar vdd precharge_0
Xpre_column_46 bl_46 br_46 en_bar vdd precharge_0
Xpre_column_47 bl_47 br_47 en_bar vdd precharge_0
Xpre_column_48 bl_48 br_48 en_bar vdd precharge_0
Xpre_column_49 bl_49 br_49 en_bar vdd precharge_0
Xpre_column_50 bl_50 br_50 en_bar vdd precharge_0
Xpre_column_51 bl_51 br_51 en_bar vdd precharge_0
Xpre_column_52 bl_52 br_52 en_bar vdd precharge_0
Xpre_column_53 bl_53 br_53 en_bar vdd precharge_0
Xpre_column_54 bl_54 br_54 en_bar vdd precharge_0
Xpre_column_55 bl_55 br_55 en_bar vdd precharge_0
Xpre_column_56 bl_56 br_56 en_bar vdd precharge_0
Xpre_column_57 bl_57 br_57 en_bar vdd precharge_0
Xpre_column_58 bl_58 br_58 en_bar vdd precharge_0
Xpre_column_59 bl_59 br_59 en_bar vdd precharge_0
Xpre_column_60 bl_60 br_60 en_bar vdd precharge_0
Xpre_column_61 bl_61 br_61 en_bar vdd precharge_0
Xpre_column_62 bl_62 br_62 en_bar vdd precharge_0
Xpre_column_63 bl_63 br_63 en_bar vdd precharge_0
Xpre_column_64 bl_64 br_64 en_bar vdd precharge_0
Xpre_column_65 bl_65 br_65 en_bar vdd precharge_0
Xpre_column_66 bl_66 br_66 en_bar vdd precharge_0
Xpre_column_67 bl_67 br_67 en_bar vdd precharge_0
Xpre_column_68 bl_68 br_68 en_bar vdd precharge_0
Xpre_column_69 bl_69 br_69 en_bar vdd precharge_0
Xpre_column_70 bl_70 br_70 en_bar vdd precharge_0
Xpre_column_71 bl_71 br_71 en_bar vdd precharge_0
Xpre_column_72 bl_72 br_72 en_bar vdd precharge_0
Xpre_column_73 bl_73 br_73 en_bar vdd precharge_0
Xpre_column_74 bl_74 br_74 en_bar vdd precharge_0
Xpre_column_75 bl_75 br_75 en_bar vdd precharge_0
Xpre_column_76 bl_76 br_76 en_bar vdd precharge_0
Xpre_column_77 bl_77 br_77 en_bar vdd precharge_0
Xpre_column_78 bl_78 br_78 en_bar vdd precharge_0
Xpre_column_79 bl_79 br_79 en_bar vdd precharge_0
Xpre_column_80 bl_80 br_80 en_bar vdd precharge_0
Xpre_column_81 bl_81 br_81 en_bar vdd precharge_0
Xpre_column_82 bl_82 br_82 en_bar vdd precharge_0
Xpre_column_83 bl_83 br_83 en_bar vdd precharge_0
Xpre_column_84 bl_84 br_84 en_bar vdd precharge_0
Xpre_column_85 bl_85 br_85 en_bar vdd precharge_0
Xpre_column_86 bl_86 br_86 en_bar vdd precharge_0
Xpre_column_87 bl_87 br_87 en_bar vdd precharge_0
Xpre_column_88 bl_88 br_88 en_bar vdd precharge_0
Xpre_column_89 bl_89 br_89 en_bar vdd precharge_0
Xpre_column_90 bl_90 br_90 en_bar vdd precharge_0
Xpre_column_91 bl_91 br_91 en_bar vdd precharge_0
Xpre_column_92 bl_92 br_92 en_bar vdd precharge_0
Xpre_column_93 bl_93 br_93 en_bar vdd precharge_0
Xpre_column_94 bl_94 br_94 en_bar vdd precharge_0
Xpre_column_95 bl_95 br_95 en_bar vdd precharge_0
Xpre_column_96 bl_96 br_96 en_bar vdd precharge_0
Xpre_column_97 bl_97 br_97 en_bar vdd precharge_0
Xpre_column_98 bl_98 br_98 en_bar vdd precharge_0
Xpre_column_99 bl_99 br_99 en_bar vdd precharge_0
Xpre_column_100 bl_100 br_100 en_bar vdd precharge_0
Xpre_column_101 bl_101 br_101 en_bar vdd precharge_0
Xpre_column_102 bl_102 br_102 en_bar vdd precharge_0
Xpre_column_103 bl_103 br_103 en_bar vdd precharge_0
Xpre_column_104 bl_104 br_104 en_bar vdd precharge_0
Xpre_column_105 bl_105 br_105 en_bar vdd precharge_0
Xpre_column_106 bl_106 br_106 en_bar vdd precharge_0
Xpre_column_107 bl_107 br_107 en_bar vdd precharge_0
Xpre_column_108 bl_108 br_108 en_bar vdd precharge_0
Xpre_column_109 bl_109 br_109 en_bar vdd precharge_0
Xpre_column_110 bl_110 br_110 en_bar vdd precharge_0
Xpre_column_111 bl_111 br_111 en_bar vdd precharge_0
Xpre_column_112 bl_112 br_112 en_bar vdd precharge_0
Xpre_column_113 bl_113 br_113 en_bar vdd precharge_0
Xpre_column_114 bl_114 br_114 en_bar vdd precharge_0
Xpre_column_115 bl_115 br_115 en_bar vdd precharge_0
Xpre_column_116 bl_116 br_116 en_bar vdd precharge_0
Xpre_column_117 bl_117 br_117 en_bar vdd precharge_0
Xpre_column_118 bl_118 br_118 en_bar vdd precharge_0
Xpre_column_119 bl_119 br_119 en_bar vdd precharge_0
Xpre_column_120 bl_120 br_120 en_bar vdd precharge_0
Xpre_column_121 bl_121 br_121 en_bar vdd precharge_0
Xpre_column_122 bl_122 br_122 en_bar vdd precharge_0
Xpre_column_123 bl_123 br_123 en_bar vdd precharge_0
Xpre_column_124 bl_124 br_124 en_bar vdd precharge_0
Xpre_column_125 bl_125 br_125 en_bar vdd precharge_0
Xpre_column_126 bl_126 br_126 en_bar vdd precharge_0
Xpre_column_127 bl_127 br_127 en_bar vdd precharge_0
Xpre_column_128 bl_128 br_128 en_bar vdd precharge_0
Xpre_column_129 bl_129 br_129 en_bar vdd precharge_0
.ENDS precharge_array
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

*********************** "sky130_fd_bd_sram__openram_sense_amp" ******************************

.SUBCKT sky130_fd_bd_sram__openram_sense_amp BL BR DOUT EN VDD GND
X1000 GND EN a_56_432# GND sky130_fd_pr__nfet_01v8 W=0.65 L=0.15
X1001 a_56_432# dint_bar dint GND sky130_fd_pr__nfet_01v8 W=0.65 L=0.15
X1002 dint_bar dint a_56_432# GND sky130_fd_pr__nfet_01v8 W=0.65 L=0.15

X1003 VDD dint_bar dint VDD sky130_fd_pr__pfet_01v8 W=1.26 L=0.15
X1004 dint_bar dint VDD VDD sky130_fd_pr__pfet_01v8 W=1.26 L=0.15

X1005 BL EN dint VDD sky130_fd_pr__pfet_01v8 W=2 L=0.15
X1006 dint_bar EN BR VDD sky130_fd_pr__pfet_01v8 W=2 L=0.15

X1007 VDD dint_bar DOUT VDD sky130_fd_pr__pfet_01v8 W=1.26 L=0.15
X1008 DOUT dint_bar GND GND sky130_fd_pr__nfet_01v8 W=0.65 L=0.15

.ENDS sky130_fd_bd_sram__openram_sense_amp

.SUBCKT sense_amp_array data_0 bl_0 br_0 data_1 bl_1 br_1 data_2 bl_2 br_2 data_3 bl_3 br_3 data_4 bl_4 br_4 data_5 bl_5 br_5 data_6 bl_6 br_6 data_7 bl_7 br_7 data_8 bl_8 br_8 data_9 bl_9 br_9 data_10 bl_10 br_10 data_11 bl_11 br_11 data_12 bl_12 br_12 data_13 bl_13 br_13 data_14 bl_14 br_14 data_15 bl_15 br_15 data_16 bl_16 br_16 data_17 bl_17 br_17 data_18 bl_18 br_18 data_19 bl_19 br_19 data_20 bl_20 br_20 data_21 bl_21 br_21 data_22 bl_22 br_22 data_23 bl_23 br_23 data_24 bl_24 br_24 data_25 bl_25 br_25 data_26 bl_26 br_26 data_27 bl_27 br_27 data_28 bl_28 br_28 data_29 bl_29 br_29 data_30 bl_30 br_30 data_31 bl_31 br_31 data_32 bl_32 br_32 en vdd gnd
*.PININFO data_0:O bl_0:I br_0:I data_1:O bl_1:I br_1:I data_2:O bl_2:I br_2:I data_3:O bl_3:I br_3:I data_4:O bl_4:I br_4:I data_5:O bl_5:I br_5:I data_6:O bl_6:I br_6:I data_7:O bl_7:I br_7:I data_8:O bl_8:I br_8:I data_9:O bl_9:I br_9:I data_10:O bl_10:I br_10:I data_11:O bl_11:I br_11:I data_12:O bl_12:I br_12:I data_13:O bl_13:I br_13:I data_14:O bl_14:I br_14:I data_15:O bl_15:I br_15:I data_16:O bl_16:I br_16:I data_17:O bl_17:I br_17:I data_18:O bl_18:I br_18:I data_19:O bl_19:I br_19:I data_20:O bl_20:I br_20:I data_21:O bl_21:I br_21:I data_22:O bl_22:I br_22:I data_23:O bl_23:I br_23:I data_24:O bl_24:I br_24:I data_25:O bl_25:I br_25:I data_26:O bl_26:I br_26:I data_27:O bl_27:I br_27:I data_28:O bl_28:I br_28:I data_29:O bl_29:I br_29:I data_30:O bl_30:I br_30:I data_31:O bl_31:I br_31:I data_32:O bl_32:I br_32:I en:I vdd:B gnd:B
* OUTPUT: data_0 
* INPUT : bl_0 
* INPUT : br_0 
* OUTPUT: data_1 
* INPUT : bl_1 
* INPUT : br_1 
* OUTPUT: data_2 
* INPUT : bl_2 
* INPUT : br_2 
* OUTPUT: data_3 
* INPUT : bl_3 
* INPUT : br_3 
* OUTPUT: data_4 
* INPUT : bl_4 
* INPUT : br_4 
* OUTPUT: data_5 
* INPUT : bl_5 
* INPUT : br_5 
* OUTPUT: data_6 
* INPUT : bl_6 
* INPUT : br_6 
* OUTPUT: data_7 
* INPUT : bl_7 
* INPUT : br_7 
* OUTPUT: data_8 
* INPUT : bl_8 
* INPUT : br_8 
* OUTPUT: data_9 
* INPUT : bl_9 
* INPUT : br_9 
* OUTPUT: data_10 
* INPUT : bl_10 
* INPUT : br_10 
* OUTPUT: data_11 
* INPUT : bl_11 
* INPUT : br_11 
* OUTPUT: data_12 
* INPUT : bl_12 
* INPUT : br_12 
* OUTPUT: data_13 
* INPUT : bl_13 
* INPUT : br_13 
* OUTPUT: data_14 
* INPUT : bl_14 
* INPUT : br_14 
* OUTPUT: data_15 
* INPUT : bl_15 
* INPUT : br_15 
* OUTPUT: data_16 
* INPUT : bl_16 
* INPUT : br_16 
* OUTPUT: data_17 
* INPUT : bl_17 
* INPUT : br_17 
* OUTPUT: data_18 
* INPUT : bl_18 
* INPUT : br_18 
* OUTPUT: data_19 
* INPUT : bl_19 
* INPUT : br_19 
* OUTPUT: data_20 
* INPUT : bl_20 
* INPUT : br_20 
* OUTPUT: data_21 
* INPUT : bl_21 
* INPUT : br_21 
* OUTPUT: data_22 
* INPUT : bl_22 
* INPUT : br_22 
* OUTPUT: data_23 
* INPUT : bl_23 
* INPUT : br_23 
* OUTPUT: data_24 
* INPUT : bl_24 
* INPUT : br_24 
* OUTPUT: data_25 
* INPUT : bl_25 
* INPUT : br_25 
* OUTPUT: data_26 
* INPUT : bl_26 
* INPUT : br_26 
* OUTPUT: data_27 
* INPUT : bl_27 
* INPUT : br_27 
* OUTPUT: data_28 
* INPUT : bl_28 
* INPUT : br_28 
* OUTPUT: data_29 
* INPUT : bl_29 
* INPUT : br_29 
* OUTPUT: data_30 
* INPUT : bl_30 
* INPUT : br_30 
* OUTPUT: data_31 
* INPUT : bl_31 
* INPUT : br_31 
* OUTPUT: data_32 
* INPUT : bl_32 
* INPUT : br_32 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* words_per_row: 4
Xsa_d0 bl_0 br_0 data_0 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d1 bl_1 br_1 data_1 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d2 bl_2 br_2 data_2 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d3 bl_3 br_3 data_3 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d4 bl_4 br_4 data_4 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d5 bl_5 br_5 data_5 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d6 bl_6 br_6 data_6 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d7 bl_7 br_7 data_7 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d8 bl_8 br_8 data_8 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d9 bl_9 br_9 data_9 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d10 bl_10 br_10 data_10 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d11 bl_11 br_11 data_11 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d12 bl_12 br_12 data_12 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d13 bl_13 br_13 data_13 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d14 bl_14 br_14 data_14 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d15 bl_15 br_15 data_15 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d16 bl_16 br_16 data_16 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d17 bl_17 br_17 data_17 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d18 bl_18 br_18 data_18 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d19 bl_19 br_19 data_19 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d20 bl_20 br_20 data_20 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d21 bl_21 br_21 data_21 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d22 bl_22 br_22 data_22 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d23 bl_23 br_23 data_23 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d24 bl_24 br_24 data_24 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d25 bl_25 br_25 data_25 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d26 bl_26 br_26 data_26 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d27 bl_27 br_27 data_27 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d28 bl_28 br_28 data_28 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d29 bl_29 br_29 data_29 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d30 bl_30 br_30 data_30 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d31 bl_31 br_31 data_31 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsa_d32 bl_32 br_32 data_32 en vdd gnd sky130_fd_bd_sram__openram_sense_amp
.ENDS sense_amp_array

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.88 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u

.SUBCKT column_mux bl br bl_out br_out sel gnd
*.PININFO bl:B br:B bl_out:B br_out:B sel:B gnd:B
* INOUT : bl 
* INOUT : br 
* INOUT : bl_out 
* INOUT : br_out 
* INOUT : sel 
* INOUT : gnd 
Xmux_tx1 bl sel bl_out gnd sky130_fd_pr__nfet_01v8 m=1 w=2.88 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u
Xmux_tx2 br sel br_out gnd sky130_fd_pr__nfet_01v8 m=1 w=2.88 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u
.ENDS column_mux

.SUBCKT column_mux_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 sel_0 sel_1 sel_2 sel_3 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 gnd
*.PININFO bl_0:B br_0:B bl_1:B br_1:B bl_2:B br_2:B bl_3:B br_3:B bl_4:B br_4:B bl_5:B br_5:B bl_6:B br_6:B bl_7:B br_7:B bl_8:B br_8:B bl_9:B br_9:B bl_10:B br_10:B bl_11:B br_11:B bl_12:B br_12:B bl_13:B br_13:B bl_14:B br_14:B bl_15:B br_15:B bl_16:B br_16:B bl_17:B br_17:B bl_18:B br_18:B bl_19:B br_19:B bl_20:B br_20:B bl_21:B br_21:B bl_22:B br_22:B bl_23:B br_23:B bl_24:B br_24:B bl_25:B br_25:B bl_26:B br_26:B bl_27:B br_27:B bl_28:B br_28:B bl_29:B br_29:B bl_30:B br_30:B bl_31:B br_31:B bl_32:B br_32:B bl_33:B br_33:B bl_34:B br_34:B bl_35:B br_35:B bl_36:B br_36:B bl_37:B br_37:B bl_38:B br_38:B bl_39:B br_39:B bl_40:B br_40:B bl_41:B br_41:B bl_42:B br_42:B bl_43:B br_43:B bl_44:B br_44:B bl_45:B br_45:B bl_46:B br_46:B bl_47:B br_47:B bl_48:B br_48:B bl_49:B br_49:B bl_50:B br_50:B bl_51:B br_51:B bl_52:B br_52:B bl_53:B br_53:B bl_54:B br_54:B bl_55:B br_55:B bl_56:B br_56:B bl_57:B br_57:B bl_58:B br_58:B bl_59:B br_59:B bl_60:B br_60:B bl_61:B br_61:B bl_62:B br_62:B bl_63:B br_63:B bl_64:B br_64:B bl_65:B br_65:B bl_66:B br_66:B bl_67:B br_67:B bl_68:B br_68:B bl_69:B br_69:B bl_70:B br_70:B bl_71:B br_71:B bl_72:B br_72:B bl_73:B br_73:B bl_74:B br_74:B bl_75:B br_75:B bl_76:B br_76:B bl_77:B br_77:B bl_78:B br_78:B bl_79:B br_79:B bl_80:B br_80:B bl_81:B br_81:B bl_82:B br_82:B bl_83:B br_83:B bl_84:B br_84:B bl_85:B br_85:B bl_86:B br_86:B bl_87:B br_87:B bl_88:B br_88:B bl_89:B br_89:B bl_90:B br_90:B bl_91:B br_91:B bl_92:B br_92:B bl_93:B br_93:B bl_94:B br_94:B bl_95:B br_95:B bl_96:B br_96:B bl_97:B br_97:B bl_98:B br_98:B bl_99:B br_99:B bl_100:B br_100:B bl_101:B br_101:B bl_102:B br_102:B bl_103:B br_103:B bl_104:B br_104:B bl_105:B br_105:B bl_106:B br_106:B bl_107:B br_107:B bl_108:B br_108:B bl_109:B br_109:B bl_110:B br_110:B bl_111:B br_111:B bl_112:B br_112:B bl_113:B br_113:B bl_114:B br_114:B bl_115:B br_115:B bl_116:B br_116:B bl_117:B br_117:B bl_118:B br_118:B bl_119:B br_119:B bl_120:B br_120:B bl_121:B br_121:B bl_122:B br_122:B bl_123:B br_123:B bl_124:B br_124:B bl_125:B br_125:B bl_126:B br_126:B bl_127:B br_127:B sel_0:B sel_1:B sel_2:B sel_3:B bl_out_0:B br_out_0:B bl_out_1:B br_out_1:B bl_out_2:B br_out_2:B bl_out_3:B br_out_3:B bl_out_4:B br_out_4:B bl_out_5:B br_out_5:B bl_out_6:B br_out_6:B bl_out_7:B br_out_7:B bl_out_8:B br_out_8:B bl_out_9:B br_out_9:B bl_out_10:B br_out_10:B bl_out_11:B br_out_11:B bl_out_12:B br_out_12:B bl_out_13:B br_out_13:B bl_out_14:B br_out_14:B bl_out_15:B br_out_15:B bl_out_16:B br_out_16:B bl_out_17:B br_out_17:B bl_out_18:B br_out_18:B bl_out_19:B br_out_19:B bl_out_20:B br_out_20:B bl_out_21:B br_out_21:B bl_out_22:B br_out_22:B bl_out_23:B br_out_23:B bl_out_24:B br_out_24:B bl_out_25:B br_out_25:B bl_out_26:B br_out_26:B bl_out_27:B br_out_27:B bl_out_28:B br_out_28:B bl_out_29:B br_out_29:B bl_out_30:B br_out_30:B bl_out_31:B br_out_31:B gnd:B
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : sel_0 
* INOUT : sel_1 
* INOUT : sel_2 
* INOUT : sel_3 
* INOUT : bl_out_0 
* INOUT : br_out_0 
* INOUT : bl_out_1 
* INOUT : br_out_1 
* INOUT : bl_out_2 
* INOUT : br_out_2 
* INOUT : bl_out_3 
* INOUT : br_out_3 
* INOUT : bl_out_4 
* INOUT : br_out_4 
* INOUT : bl_out_5 
* INOUT : br_out_5 
* INOUT : bl_out_6 
* INOUT : br_out_6 
* INOUT : bl_out_7 
* INOUT : br_out_7 
* INOUT : bl_out_8 
* INOUT : br_out_8 
* INOUT : bl_out_9 
* INOUT : br_out_9 
* INOUT : bl_out_10 
* INOUT : br_out_10 
* INOUT : bl_out_11 
* INOUT : br_out_11 
* INOUT : bl_out_12 
* INOUT : br_out_12 
* INOUT : bl_out_13 
* INOUT : br_out_13 
* INOUT : bl_out_14 
* INOUT : br_out_14 
* INOUT : bl_out_15 
* INOUT : br_out_15 
* INOUT : bl_out_16 
* INOUT : br_out_16 
* INOUT : bl_out_17 
* INOUT : br_out_17 
* INOUT : bl_out_18 
* INOUT : br_out_18 
* INOUT : bl_out_19 
* INOUT : br_out_19 
* INOUT : bl_out_20 
* INOUT : br_out_20 
* INOUT : bl_out_21 
* INOUT : br_out_21 
* INOUT : bl_out_22 
* INOUT : br_out_22 
* INOUT : bl_out_23 
* INOUT : br_out_23 
* INOUT : bl_out_24 
* INOUT : br_out_24 
* INOUT : bl_out_25 
* INOUT : br_out_25 
* INOUT : bl_out_26 
* INOUT : br_out_26 
* INOUT : bl_out_27 
* INOUT : br_out_27 
* INOUT : bl_out_28 
* INOUT : br_out_28 
* INOUT : bl_out_29 
* INOUT : br_out_29 
* INOUT : bl_out_30 
* INOUT : br_out_30 
* INOUT : bl_out_31 
* INOUT : br_out_31 
* INOUT : gnd 
* cols: 128 word_size: 32 bl: bl br: br
XXMUX0 bl_0 br_0 bl_out_0 br_out_0 sel_0 gnd column_mux
XXMUX1 bl_1 br_1 bl_out_0 br_out_0 sel_1 gnd column_mux
XXMUX2 bl_2 br_2 bl_out_0 br_out_0 sel_2 gnd column_mux
XXMUX3 bl_3 br_3 bl_out_0 br_out_0 sel_3 gnd column_mux
XXMUX4 bl_4 br_4 bl_out_1 br_out_1 sel_0 gnd column_mux
XXMUX5 bl_5 br_5 bl_out_1 br_out_1 sel_1 gnd column_mux
XXMUX6 bl_6 br_6 bl_out_1 br_out_1 sel_2 gnd column_mux
XXMUX7 bl_7 br_7 bl_out_1 br_out_1 sel_3 gnd column_mux
XXMUX8 bl_8 br_8 bl_out_2 br_out_2 sel_0 gnd column_mux
XXMUX9 bl_9 br_9 bl_out_2 br_out_2 sel_1 gnd column_mux
XXMUX10 bl_10 br_10 bl_out_2 br_out_2 sel_2 gnd column_mux
XXMUX11 bl_11 br_11 bl_out_2 br_out_2 sel_3 gnd column_mux
XXMUX12 bl_12 br_12 bl_out_3 br_out_3 sel_0 gnd column_mux
XXMUX13 bl_13 br_13 bl_out_3 br_out_3 sel_1 gnd column_mux
XXMUX14 bl_14 br_14 bl_out_3 br_out_3 sel_2 gnd column_mux
XXMUX15 bl_15 br_15 bl_out_3 br_out_3 sel_3 gnd column_mux
XXMUX16 bl_16 br_16 bl_out_4 br_out_4 sel_0 gnd column_mux
XXMUX17 bl_17 br_17 bl_out_4 br_out_4 sel_1 gnd column_mux
XXMUX18 bl_18 br_18 bl_out_4 br_out_4 sel_2 gnd column_mux
XXMUX19 bl_19 br_19 bl_out_4 br_out_4 sel_3 gnd column_mux
XXMUX20 bl_20 br_20 bl_out_5 br_out_5 sel_0 gnd column_mux
XXMUX21 bl_21 br_21 bl_out_5 br_out_5 sel_1 gnd column_mux
XXMUX22 bl_22 br_22 bl_out_5 br_out_5 sel_2 gnd column_mux
XXMUX23 bl_23 br_23 bl_out_5 br_out_5 sel_3 gnd column_mux
XXMUX24 bl_24 br_24 bl_out_6 br_out_6 sel_0 gnd column_mux
XXMUX25 bl_25 br_25 bl_out_6 br_out_6 sel_1 gnd column_mux
XXMUX26 bl_26 br_26 bl_out_6 br_out_6 sel_2 gnd column_mux
XXMUX27 bl_27 br_27 bl_out_6 br_out_6 sel_3 gnd column_mux
XXMUX28 bl_28 br_28 bl_out_7 br_out_7 sel_0 gnd column_mux
XXMUX29 bl_29 br_29 bl_out_7 br_out_7 sel_1 gnd column_mux
XXMUX30 bl_30 br_30 bl_out_7 br_out_7 sel_2 gnd column_mux
XXMUX31 bl_31 br_31 bl_out_7 br_out_7 sel_3 gnd column_mux
XXMUX32 bl_32 br_32 bl_out_8 br_out_8 sel_0 gnd column_mux
XXMUX33 bl_33 br_33 bl_out_8 br_out_8 sel_1 gnd column_mux
XXMUX34 bl_34 br_34 bl_out_8 br_out_8 sel_2 gnd column_mux
XXMUX35 bl_35 br_35 bl_out_8 br_out_8 sel_3 gnd column_mux
XXMUX36 bl_36 br_36 bl_out_9 br_out_9 sel_0 gnd column_mux
XXMUX37 bl_37 br_37 bl_out_9 br_out_9 sel_1 gnd column_mux
XXMUX38 bl_38 br_38 bl_out_9 br_out_9 sel_2 gnd column_mux
XXMUX39 bl_39 br_39 bl_out_9 br_out_9 sel_3 gnd column_mux
XXMUX40 bl_40 br_40 bl_out_10 br_out_10 sel_0 gnd column_mux
XXMUX41 bl_41 br_41 bl_out_10 br_out_10 sel_1 gnd column_mux
XXMUX42 bl_42 br_42 bl_out_10 br_out_10 sel_2 gnd column_mux
XXMUX43 bl_43 br_43 bl_out_10 br_out_10 sel_3 gnd column_mux
XXMUX44 bl_44 br_44 bl_out_11 br_out_11 sel_0 gnd column_mux
XXMUX45 bl_45 br_45 bl_out_11 br_out_11 sel_1 gnd column_mux
XXMUX46 bl_46 br_46 bl_out_11 br_out_11 sel_2 gnd column_mux
XXMUX47 bl_47 br_47 bl_out_11 br_out_11 sel_3 gnd column_mux
XXMUX48 bl_48 br_48 bl_out_12 br_out_12 sel_0 gnd column_mux
XXMUX49 bl_49 br_49 bl_out_12 br_out_12 sel_1 gnd column_mux
XXMUX50 bl_50 br_50 bl_out_12 br_out_12 sel_2 gnd column_mux
XXMUX51 bl_51 br_51 bl_out_12 br_out_12 sel_3 gnd column_mux
XXMUX52 bl_52 br_52 bl_out_13 br_out_13 sel_0 gnd column_mux
XXMUX53 bl_53 br_53 bl_out_13 br_out_13 sel_1 gnd column_mux
XXMUX54 bl_54 br_54 bl_out_13 br_out_13 sel_2 gnd column_mux
XXMUX55 bl_55 br_55 bl_out_13 br_out_13 sel_3 gnd column_mux
XXMUX56 bl_56 br_56 bl_out_14 br_out_14 sel_0 gnd column_mux
XXMUX57 bl_57 br_57 bl_out_14 br_out_14 sel_1 gnd column_mux
XXMUX58 bl_58 br_58 bl_out_14 br_out_14 sel_2 gnd column_mux
XXMUX59 bl_59 br_59 bl_out_14 br_out_14 sel_3 gnd column_mux
XXMUX60 bl_60 br_60 bl_out_15 br_out_15 sel_0 gnd column_mux
XXMUX61 bl_61 br_61 bl_out_15 br_out_15 sel_1 gnd column_mux
XXMUX62 bl_62 br_62 bl_out_15 br_out_15 sel_2 gnd column_mux
XXMUX63 bl_63 br_63 bl_out_15 br_out_15 sel_3 gnd column_mux
XXMUX64 bl_64 br_64 bl_out_16 br_out_16 sel_0 gnd column_mux
XXMUX65 bl_65 br_65 bl_out_16 br_out_16 sel_1 gnd column_mux
XXMUX66 bl_66 br_66 bl_out_16 br_out_16 sel_2 gnd column_mux
XXMUX67 bl_67 br_67 bl_out_16 br_out_16 sel_3 gnd column_mux
XXMUX68 bl_68 br_68 bl_out_17 br_out_17 sel_0 gnd column_mux
XXMUX69 bl_69 br_69 bl_out_17 br_out_17 sel_1 gnd column_mux
XXMUX70 bl_70 br_70 bl_out_17 br_out_17 sel_2 gnd column_mux
XXMUX71 bl_71 br_71 bl_out_17 br_out_17 sel_3 gnd column_mux
XXMUX72 bl_72 br_72 bl_out_18 br_out_18 sel_0 gnd column_mux
XXMUX73 bl_73 br_73 bl_out_18 br_out_18 sel_1 gnd column_mux
XXMUX74 bl_74 br_74 bl_out_18 br_out_18 sel_2 gnd column_mux
XXMUX75 bl_75 br_75 bl_out_18 br_out_18 sel_3 gnd column_mux
XXMUX76 bl_76 br_76 bl_out_19 br_out_19 sel_0 gnd column_mux
XXMUX77 bl_77 br_77 bl_out_19 br_out_19 sel_1 gnd column_mux
XXMUX78 bl_78 br_78 bl_out_19 br_out_19 sel_2 gnd column_mux
XXMUX79 bl_79 br_79 bl_out_19 br_out_19 sel_3 gnd column_mux
XXMUX80 bl_80 br_80 bl_out_20 br_out_20 sel_0 gnd column_mux
XXMUX81 bl_81 br_81 bl_out_20 br_out_20 sel_1 gnd column_mux
XXMUX82 bl_82 br_82 bl_out_20 br_out_20 sel_2 gnd column_mux
XXMUX83 bl_83 br_83 bl_out_20 br_out_20 sel_3 gnd column_mux
XXMUX84 bl_84 br_84 bl_out_21 br_out_21 sel_0 gnd column_mux
XXMUX85 bl_85 br_85 bl_out_21 br_out_21 sel_1 gnd column_mux
XXMUX86 bl_86 br_86 bl_out_21 br_out_21 sel_2 gnd column_mux
XXMUX87 bl_87 br_87 bl_out_21 br_out_21 sel_3 gnd column_mux
XXMUX88 bl_88 br_88 bl_out_22 br_out_22 sel_0 gnd column_mux
XXMUX89 bl_89 br_89 bl_out_22 br_out_22 sel_1 gnd column_mux
XXMUX90 bl_90 br_90 bl_out_22 br_out_22 sel_2 gnd column_mux
XXMUX91 bl_91 br_91 bl_out_22 br_out_22 sel_3 gnd column_mux
XXMUX92 bl_92 br_92 bl_out_23 br_out_23 sel_0 gnd column_mux
XXMUX93 bl_93 br_93 bl_out_23 br_out_23 sel_1 gnd column_mux
XXMUX94 bl_94 br_94 bl_out_23 br_out_23 sel_2 gnd column_mux
XXMUX95 bl_95 br_95 bl_out_23 br_out_23 sel_3 gnd column_mux
XXMUX96 bl_96 br_96 bl_out_24 br_out_24 sel_0 gnd column_mux
XXMUX97 bl_97 br_97 bl_out_24 br_out_24 sel_1 gnd column_mux
XXMUX98 bl_98 br_98 bl_out_24 br_out_24 sel_2 gnd column_mux
XXMUX99 bl_99 br_99 bl_out_24 br_out_24 sel_3 gnd column_mux
XXMUX100 bl_100 br_100 bl_out_25 br_out_25 sel_0 gnd column_mux
XXMUX101 bl_101 br_101 bl_out_25 br_out_25 sel_1 gnd column_mux
XXMUX102 bl_102 br_102 bl_out_25 br_out_25 sel_2 gnd column_mux
XXMUX103 bl_103 br_103 bl_out_25 br_out_25 sel_3 gnd column_mux
XXMUX104 bl_104 br_104 bl_out_26 br_out_26 sel_0 gnd column_mux
XXMUX105 bl_105 br_105 bl_out_26 br_out_26 sel_1 gnd column_mux
XXMUX106 bl_106 br_106 bl_out_26 br_out_26 sel_2 gnd column_mux
XXMUX107 bl_107 br_107 bl_out_26 br_out_26 sel_3 gnd column_mux
XXMUX108 bl_108 br_108 bl_out_27 br_out_27 sel_0 gnd column_mux
XXMUX109 bl_109 br_109 bl_out_27 br_out_27 sel_1 gnd column_mux
XXMUX110 bl_110 br_110 bl_out_27 br_out_27 sel_2 gnd column_mux
XXMUX111 bl_111 br_111 bl_out_27 br_out_27 sel_3 gnd column_mux
XXMUX112 bl_112 br_112 bl_out_28 br_out_28 sel_0 gnd column_mux
XXMUX113 bl_113 br_113 bl_out_28 br_out_28 sel_1 gnd column_mux
XXMUX114 bl_114 br_114 bl_out_28 br_out_28 sel_2 gnd column_mux
XXMUX115 bl_115 br_115 bl_out_28 br_out_28 sel_3 gnd column_mux
XXMUX116 bl_116 br_116 bl_out_29 br_out_29 sel_0 gnd column_mux
XXMUX117 bl_117 br_117 bl_out_29 br_out_29 sel_1 gnd column_mux
XXMUX118 bl_118 br_118 bl_out_29 br_out_29 sel_2 gnd column_mux
XXMUX119 bl_119 br_119 bl_out_29 br_out_29 sel_3 gnd column_mux
XXMUX120 bl_120 br_120 bl_out_30 br_out_30 sel_0 gnd column_mux
XXMUX121 bl_121 br_121 bl_out_30 br_out_30 sel_1 gnd column_mux
XXMUX122 bl_122 br_122 bl_out_30 br_out_30 sel_2 gnd column_mux
XXMUX123 bl_123 br_123 bl_out_30 br_out_30 sel_3 gnd column_mux
XXMUX124 bl_124 br_124 bl_out_31 br_out_31 sel_0 gnd column_mux
XXMUX125 bl_125 br_125 bl_out_31 br_out_31 sel_1 gnd column_mux
XXMUX126 bl_126 br_126 bl_out_31 br_out_31 sel_2 gnd column_mux
XXMUX127 bl_127 br_127 bl_out_31 br_out_31 sel_3 gnd column_mux
.ENDS column_mux_array
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

*********************** "sky130_fd_bd_sram__openram_write_driver" ******************************

.SUBCKT sky130_fd_bd_sram__openram_write_driver DIN BL BR EN VDD GND

**** Inverter to conver Data_in to data_in_bar ******
* din_bar = inv(DIN)
X_1 din_bar DIN GND GND sky130_fd_pr__nfet_01v8 W=0.36 L=0.15
X_2 din_bar DIN VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15

**** 2input nand gate follwed by inverter to drive BL ******
* din_bar_gated = nand(EN, DIN)
X_3 din_bar_gated EN net_7 GND sky130_fd_pr__nfet_01v8 W=0.55 L=0.15
X_4 net_7 DIN GND GND sky130_fd_pr__nfet_01v8 W=0.55 L=0.15
X_5 din_bar_gated EN VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
X_6 din_bar_gated DIN VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
* din_bar_gated_bar = inv(din_bar_gated)
X_7 din_bar_gated_bar din_bar_gated VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
X_8 din_bar_gated_bar din_bar_gated GND GND sky130_fd_pr__nfet_01v8 W=0.36 L=0.15

**** 2input nand gate follwed by inverter to drive BR******
* din_gated = nand(EN, din_bar)
X_9 din_gated EN VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
X_10 din_gated EN net_8 GND sky130_fd_pr__nfet_01v8 W=0.55 L=0.15
X_11 net_8 din_bar GND GND sky130_fd_pr__nfet_01v8 W=0.55 L=0.15
X_12 din_gated din_bar VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
* din_gated_bar = inv(din_gated)
X_13 din_gated_bar din_gated VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
X_14 din_gated_bar din_gated GND GND sky130_fd_pr__nfet_01v8 W=0.36 L=0.15

************************************************
* pull down with EN enable
X_15 BL din_gated_bar GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X_16 BR din_bar_gated_bar GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15

.ENDS sky130_fd_bd_sram__openram_write_driver

.SUBCKT write_driver_array data_0 data_1 data_2 data_3 data_4 data_5 data_6 data_7 data_8 data_9 data_10 data_11 data_12 data_13 data_14 data_15 data_16 data_17 data_18 data_19 data_20 data_21 data_22 data_23 data_24 data_25 data_26 data_27 data_28 data_29 data_30 data_31 data_32 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 en_0 en_1 en_2 en_3 en_4 vdd gnd
*.PININFO data_0:I data_1:I data_2:I data_3:I data_4:I data_5:I data_6:I data_7:I data_8:I data_9:I data_10:I data_11:I data_12:I data_13:I data_14:I data_15:I data_16:I data_17:I data_18:I data_19:I data_20:I data_21:I data_22:I data_23:I data_24:I data_25:I data_26:I data_27:I data_28:I data_29:I data_30:I data_31:I data_32:I bl_0:O br_0:O bl_1:O br_1:O bl_2:O br_2:O bl_3:O br_3:O bl_4:O br_4:O bl_5:O br_5:O bl_6:O br_6:O bl_7:O br_7:O bl_8:O br_8:O bl_9:O br_9:O bl_10:O br_10:O bl_11:O br_11:O bl_12:O br_12:O bl_13:O br_13:O bl_14:O br_14:O bl_15:O br_15:O bl_16:O br_16:O bl_17:O br_17:O bl_18:O br_18:O bl_19:O br_19:O bl_20:O br_20:O bl_21:O br_21:O bl_22:O br_22:O bl_23:O br_23:O bl_24:O br_24:O bl_25:O br_25:O bl_26:O br_26:O bl_27:O br_27:O bl_28:O br_28:O bl_29:O br_29:O bl_30:O br_30:O bl_31:O br_31:O bl_32:O br_32:O en_0:I en_1:I en_2:I en_3:I en_4:I vdd:B gnd:B
* INPUT : data_0 
* INPUT : data_1 
* INPUT : data_2 
* INPUT : data_3 
* INPUT : data_4 
* INPUT : data_5 
* INPUT : data_6 
* INPUT : data_7 
* INPUT : data_8 
* INPUT : data_9 
* INPUT : data_10 
* INPUT : data_11 
* INPUT : data_12 
* INPUT : data_13 
* INPUT : data_14 
* INPUT : data_15 
* INPUT : data_16 
* INPUT : data_17 
* INPUT : data_18 
* INPUT : data_19 
* INPUT : data_20 
* INPUT : data_21 
* INPUT : data_22 
* INPUT : data_23 
* INPUT : data_24 
* INPUT : data_25 
* INPUT : data_26 
* INPUT : data_27 
* INPUT : data_28 
* INPUT : data_29 
* INPUT : data_30 
* INPUT : data_31 
* INPUT : data_32 
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* INPUT : en_0 
* INPUT : en_1 
* INPUT : en_2 
* INPUT : en_3 
* INPUT : en_4 
* POWER : vdd 
* GROUND: gnd 
* word_size 32
Xwrite_driver0 data_0 bl_0 br_0 en_0 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver4 data_1 bl_1 br_1 en_0 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver8 data_2 bl_2 br_2 en_0 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver12 data_3 bl_3 br_3 en_0 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver16 data_4 bl_4 br_4 en_0 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver20 data_5 bl_5 br_5 en_0 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver24 data_6 bl_6 br_6 en_0 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver28 data_7 bl_7 br_7 en_0 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver32 data_8 bl_8 br_8 en_1 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver36 data_9 bl_9 br_9 en_1 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver40 data_10 bl_10 br_10 en_1 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver44 data_11 bl_11 br_11 en_1 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver48 data_12 bl_12 br_12 en_1 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver52 data_13 bl_13 br_13 en_1 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver56 data_14 bl_14 br_14 en_1 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver60 data_15 bl_15 br_15 en_1 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver64 data_16 bl_16 br_16 en_2 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver68 data_17 bl_17 br_17 en_2 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver72 data_18 bl_18 br_18 en_2 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver76 data_19 bl_19 br_19 en_2 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver80 data_20 bl_20 br_20 en_2 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver84 data_21 bl_21 br_21 en_2 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver88 data_22 bl_22 br_22 en_2 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver92 data_23 bl_23 br_23 en_2 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver96 data_24 bl_24 br_24 en_3 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver100 data_25 bl_25 br_25 en_3 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver104 data_26 bl_26 br_26 en_3 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver108 data_27 bl_27 br_27 en_3 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver112 data_28 bl_28 br_28 en_3 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver116 data_29 bl_29 br_29 en_3 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver120 data_30 bl_30 br_30 en_3 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver124 data_31 bl_31 br_31 en_3 vdd gnd sky130_fd_bd_sram__openram_write_driver
Xwrite_driver128 data_32 bl_32 br_32 en_4 vdd gnd sky130_fd_bd_sram__openram_write_driver
.ENDS write_driver_array

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u

.SUBCKT pnand2 A B Z vdd gnd
*.PININFO A:I B:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpnand2_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_nmos1 Z B net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand2_nmos2 net1 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pnand2

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=2 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u

.SUBCKT pinv A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=2 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pinv

.SUBCKT pdriver A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [2.0]
Xbuf_inv1 A Z vdd gnd pinv
.ENDS pdriver

.SUBCKT pand2 A B Z vdd gnd
*.PININFO A:I B:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand2_nand A B zb_int vdd gnd pnand2
Xpand2_inv zb_int Z vdd gnd pdriver
.ENDS pand2

.SUBCKT write_mask_and_array wmask_in_0 wmask_in_1 wmask_in_2 wmask_in_3 en wmask_out_0 wmask_out_1 wmask_out_2 wmask_out_3 vdd gnd
*.PININFO wmask_in_0:I wmask_in_1:I wmask_in_2:I wmask_in_3:I en:I wmask_out_0:O wmask_out_1:O wmask_out_2:O wmask_out_3:O vdd:B gnd:B
* INPUT : wmask_in_0 
* INPUT : wmask_in_1 
* INPUT : wmask_in_2 
* INPUT : wmask_in_3 
* INPUT : en 
* OUTPUT: wmask_out_0 
* OUTPUT: wmask_out_1 
* OUTPUT: wmask_out_2 
* OUTPUT: wmask_out_3 
* POWER : vdd 
* GROUND: gnd 
* write_size 8
Xand2_0 wmask_in_0 en wmask_out_0 vdd gnd pand2
Xand2_1 wmask_in_1 en wmask_out_1 vdd gnd pand2
Xand2_2 wmask_in_2 en wmask_out_2 vdd gnd pand2
Xand2_3 wmask_in_3 en wmask_out_3 vdd gnd pand2
.ENDS write_mask_and_array

.SUBCKT port_data rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 sparebl_0 sparebr_0 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 dout_32 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 din_32 sel_0 sel_1 sel_2 sel_3 s_en p_en_bar w_en bank_wmask_0 bank_wmask_1 bank_wmask_2 bank_wmask_3 bank_spare_wen0 vdd gnd
*.PININFO rbl_bl:B rbl_br:B bl_0:B br_0:B bl_1:B br_1:B bl_2:B br_2:B bl_3:B br_3:B bl_4:B br_4:B bl_5:B br_5:B bl_6:B br_6:B bl_7:B br_7:B bl_8:B br_8:B bl_9:B br_9:B bl_10:B br_10:B bl_11:B br_11:B bl_12:B br_12:B bl_13:B br_13:B bl_14:B br_14:B bl_15:B br_15:B bl_16:B br_16:B bl_17:B br_17:B bl_18:B br_18:B bl_19:B br_19:B bl_20:B br_20:B bl_21:B br_21:B bl_22:B br_22:B bl_23:B br_23:B bl_24:B br_24:B bl_25:B br_25:B bl_26:B br_26:B bl_27:B br_27:B bl_28:B br_28:B bl_29:B br_29:B bl_30:B br_30:B bl_31:B br_31:B bl_32:B br_32:B bl_33:B br_33:B bl_34:B br_34:B bl_35:B br_35:B bl_36:B br_36:B bl_37:B br_37:B bl_38:B br_38:B bl_39:B br_39:B bl_40:B br_40:B bl_41:B br_41:B bl_42:B br_42:B bl_43:B br_43:B bl_44:B br_44:B bl_45:B br_45:B bl_46:B br_46:B bl_47:B br_47:B bl_48:B br_48:B bl_49:B br_49:B bl_50:B br_50:B bl_51:B br_51:B bl_52:B br_52:B bl_53:B br_53:B bl_54:B br_54:B bl_55:B br_55:B bl_56:B br_56:B bl_57:B br_57:B bl_58:B br_58:B bl_59:B br_59:B bl_60:B br_60:B bl_61:B br_61:B bl_62:B br_62:B bl_63:B br_63:B bl_64:B br_64:B bl_65:B br_65:B bl_66:B br_66:B bl_67:B br_67:B bl_68:B br_68:B bl_69:B br_69:B bl_70:B br_70:B bl_71:B br_71:B bl_72:B br_72:B bl_73:B br_73:B bl_74:B br_74:B bl_75:B br_75:B bl_76:B br_76:B bl_77:B br_77:B bl_78:B br_78:B bl_79:B br_79:B bl_80:B br_80:B bl_81:B br_81:B bl_82:B br_82:B bl_83:B br_83:B bl_84:B br_84:B bl_85:B br_85:B bl_86:B br_86:B bl_87:B br_87:B bl_88:B br_88:B bl_89:B br_89:B bl_90:B br_90:B bl_91:B br_91:B bl_92:B br_92:B bl_93:B br_93:B bl_94:B br_94:B bl_95:B br_95:B bl_96:B br_96:B bl_97:B br_97:B bl_98:B br_98:B bl_99:B br_99:B bl_100:B br_100:B bl_101:B br_101:B bl_102:B br_102:B bl_103:B br_103:B bl_104:B br_104:B bl_105:B br_105:B bl_106:B br_106:B bl_107:B br_107:B bl_108:B br_108:B bl_109:B br_109:B bl_110:B br_110:B bl_111:B br_111:B bl_112:B br_112:B bl_113:B br_113:B bl_114:B br_114:B bl_115:B br_115:B bl_116:B br_116:B bl_117:B br_117:B bl_118:B br_118:B bl_119:B br_119:B bl_120:B br_120:B bl_121:B br_121:B bl_122:B br_122:B bl_123:B br_123:B bl_124:B br_124:B bl_125:B br_125:B bl_126:B br_126:B bl_127:B br_127:B sparebl_0:B sparebr_0:B dout_0:O dout_1:O dout_2:O dout_3:O dout_4:O dout_5:O dout_6:O dout_7:O dout_8:O dout_9:O dout_10:O dout_11:O dout_12:O dout_13:O dout_14:O dout_15:O dout_16:O dout_17:O dout_18:O dout_19:O dout_20:O dout_21:O dout_22:O dout_23:O dout_24:O dout_25:O dout_26:O dout_27:O dout_28:O dout_29:O dout_30:O dout_31:O dout_32:O din_0:I din_1:I din_2:I din_3:I din_4:I din_5:I din_6:I din_7:I din_8:I din_9:I din_10:I din_11:I din_12:I din_13:I din_14:I din_15:I din_16:I din_17:I din_18:I din_19:I din_20:I din_21:I din_22:I din_23:I din_24:I din_25:I din_26:I din_27:I din_28:I din_29:I din_30:I din_31:I din_32:I sel_0:I sel_1:I sel_2:I sel_3:I s_en:I p_en_bar:I w_en:I bank_wmask_0:I bank_wmask_1:I bank_wmask_2:I bank_wmask_3:I bank_spare_wen0:I vdd:B gnd:B
* INOUT : rbl_bl 
* INOUT : rbl_br 
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : sparebl_0 
* INOUT : sparebr_0 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* OUTPUT: dout_32 
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : din_32 
* INPUT : sel_0 
* INPUT : sel_1 
* INPUT : sel_2 
* INPUT : sel_3 
* INPUT : s_en 
* INPUT : p_en_bar 
* INPUT : w_en 
* INPUT : bank_wmask_0 
* INPUT : bank_wmask_1 
* INPUT : bank_wmask_2 
* INPUT : bank_wmask_3 
* INPUT : bank_spare_wen0 
* POWER : vdd 
* GROUND: gnd 
Xprecharge_array0 rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 sparebl_0 sparebr_0 p_en_bar vdd precharge_array
Xsense_amp_array0 dout_0 bl_out_0 br_out_0 dout_1 bl_out_1 br_out_1 dout_2 bl_out_2 br_out_2 dout_3 bl_out_3 br_out_3 dout_4 bl_out_4 br_out_4 dout_5 bl_out_5 br_out_5 dout_6 bl_out_6 br_out_6 dout_7 bl_out_7 br_out_7 dout_8 bl_out_8 br_out_8 dout_9 bl_out_9 br_out_9 dout_10 bl_out_10 br_out_10 dout_11 bl_out_11 br_out_11 dout_12 bl_out_12 br_out_12 dout_13 bl_out_13 br_out_13 dout_14 bl_out_14 br_out_14 dout_15 bl_out_15 br_out_15 dout_16 bl_out_16 br_out_16 dout_17 bl_out_17 br_out_17 dout_18 bl_out_18 br_out_18 dout_19 bl_out_19 br_out_19 dout_20 bl_out_20 br_out_20 dout_21 bl_out_21 br_out_21 dout_22 bl_out_22 br_out_22 dout_23 bl_out_23 br_out_23 dout_24 bl_out_24 br_out_24 dout_25 bl_out_25 br_out_25 dout_26 bl_out_26 br_out_26 dout_27 bl_out_27 br_out_27 dout_28 bl_out_28 br_out_28 dout_29 bl_out_29 br_out_29 dout_30 bl_out_30 br_out_30 dout_31 bl_out_31 br_out_31 dout_32 sparebl_0 sparebr_0 s_en vdd gnd sense_amp_array
Xwrite_driver_array0 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 din_32 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 sparebl_0 sparebr_0 wdriver_sel_0 wdriver_sel_1 wdriver_sel_2 wdriver_sel_3 bank_spare_wen0 vdd gnd write_driver_array
Xwrite_mask_and_array0 bank_wmask_0 bank_wmask_1 bank_wmask_2 bank_wmask_3 w_en wdriver_sel_0 wdriver_sel_1 wdriver_sel_2 wdriver_sel_3 vdd gnd write_mask_and_array
Xcolumn_mux_array0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 sel_0 sel_1 sel_2 sel_3 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 gnd column_mux_array
.ENDS port_data

.SUBCKT pnand2_0 A B Z vdd gnd
*.PININFO A:I B:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpnand2_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_nmos1 Z B net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand2_nmos2 net1 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pnand2_0

.SUBCKT pinv_0 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS pinv_0

.SUBCKT pdriver_0 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1]
Xbuf_inv1 A Z vdd gnd pinv_0
.ENDS pdriver_0

.SUBCKT pand2_0 A B Z vdd gnd
*.PININFO A:I B:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand2_nand A B zb_int vdd gnd pnand2_0
Xpand2_inv zb_int Z vdd gnd pdriver_0
.ENDS pand2_0

.SUBCKT pinv_1 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS pinv_1

.SUBCKT hierarchical_predecode2x4_0 in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
*.PININFO in_0:I in_1:I out_0:O out_1:O out_2:O out_3:O vdd:B gnd:B
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_1
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_1
XXpre2x4_and_0 inbar_0 inbar_1 out_0 vdd gnd pand2_0
XXpre2x4_and_1 in_0 inbar_1 out_1 vdd gnd pand2_0
XXpre2x4_and_2 inbar_0 in_1 out_2 vdd gnd pand2_0
XXpre2x4_and_3 in_0 in_1 out_3 vdd gnd pand2_0
.ENDS hierarchical_predecode2x4_0

.SUBCKT bank dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 dout0_32 rbl_bl_0_0 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 din0_32 addr0_0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 addr0_8 addr0_9 s_en0 p_en_bar0 w_en0 bank_wmask0_0 bank_wmask0_1 bank_wmask0_2 bank_wmask0_3 bank_spare_wen0_0 wl_en0 vdd gnd
*.PININFO dout0_0:O dout0_1:O dout0_2:O dout0_3:O dout0_4:O dout0_5:O dout0_6:O dout0_7:O dout0_8:O dout0_9:O dout0_10:O dout0_11:O dout0_12:O dout0_13:O dout0_14:O dout0_15:O dout0_16:O dout0_17:O dout0_18:O dout0_19:O dout0_20:O dout0_21:O dout0_22:O dout0_23:O dout0_24:O dout0_25:O dout0_26:O dout0_27:O dout0_28:O dout0_29:O dout0_30:O dout0_31:O dout0_32:O rbl_bl_0_0:O din0_0:I din0_1:I din0_2:I din0_3:I din0_4:I din0_5:I din0_6:I din0_7:I din0_8:I din0_9:I din0_10:I din0_11:I din0_12:I din0_13:I din0_14:I din0_15:I din0_16:I din0_17:I din0_18:I din0_19:I din0_20:I din0_21:I din0_22:I din0_23:I din0_24:I din0_25:I din0_26:I din0_27:I din0_28:I din0_29:I din0_30:I din0_31:I din0_32:I addr0_0:I addr0_1:I addr0_2:I addr0_3:I addr0_4:I addr0_5:I addr0_6:I addr0_7:I addr0_8:I addr0_9:I s_en0:I p_en_bar0:I w_en0:I bank_wmask0_0:I bank_wmask0_1:I bank_wmask0_2:I bank_wmask0_3:I bank_spare_wen0_0:I wl_en0:I vdd:B gnd:B
* OUTPUT: dout0_0 
* OUTPUT: dout0_1 
* OUTPUT: dout0_2 
* OUTPUT: dout0_3 
* OUTPUT: dout0_4 
* OUTPUT: dout0_5 
* OUTPUT: dout0_6 
* OUTPUT: dout0_7 
* OUTPUT: dout0_8 
* OUTPUT: dout0_9 
* OUTPUT: dout0_10 
* OUTPUT: dout0_11 
* OUTPUT: dout0_12 
* OUTPUT: dout0_13 
* OUTPUT: dout0_14 
* OUTPUT: dout0_15 
* OUTPUT: dout0_16 
* OUTPUT: dout0_17 
* OUTPUT: dout0_18 
* OUTPUT: dout0_19 
* OUTPUT: dout0_20 
* OUTPUT: dout0_21 
* OUTPUT: dout0_22 
* OUTPUT: dout0_23 
* OUTPUT: dout0_24 
* OUTPUT: dout0_25 
* OUTPUT: dout0_26 
* OUTPUT: dout0_27 
* OUTPUT: dout0_28 
* OUTPUT: dout0_29 
* OUTPUT: dout0_30 
* OUTPUT: dout0_31 
* OUTPUT: dout0_32 
* OUTPUT: rbl_bl_0_0 
* INPUT : din0_0 
* INPUT : din0_1 
* INPUT : din0_2 
* INPUT : din0_3 
* INPUT : din0_4 
* INPUT : din0_5 
* INPUT : din0_6 
* INPUT : din0_7 
* INPUT : din0_8 
* INPUT : din0_9 
* INPUT : din0_10 
* INPUT : din0_11 
* INPUT : din0_12 
* INPUT : din0_13 
* INPUT : din0_14 
* INPUT : din0_15 
* INPUT : din0_16 
* INPUT : din0_17 
* INPUT : din0_18 
* INPUT : din0_19 
* INPUT : din0_20 
* INPUT : din0_21 
* INPUT : din0_22 
* INPUT : din0_23 
* INPUT : din0_24 
* INPUT : din0_25 
* INPUT : din0_26 
* INPUT : din0_27 
* INPUT : din0_28 
* INPUT : din0_29 
* INPUT : din0_30 
* INPUT : din0_31 
* INPUT : din0_32 
* INPUT : addr0_0 
* INPUT : addr0_1 
* INPUT : addr0_2 
* INPUT : addr0_3 
* INPUT : addr0_4 
* INPUT : addr0_5 
* INPUT : addr0_6 
* INPUT : addr0_7 
* INPUT : addr0_8 
* INPUT : addr0_9 
* INPUT : s_en0 
* INPUT : p_en_bar0 
* INPUT : w_en0 
* INPUT : bank_wmask0_0 
* INPUT : bank_wmask0_1 
* INPUT : bank_wmask0_2 
* INPUT : bank_wmask0_3 
* INPUT : bank_spare_wen0_0 
* INPUT : wl_en0 
* POWER : vdd 
* GROUND: gnd 
Xbitcell_array rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 rbl_wl0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 vdd gnd vpb vnb sky130_replica_bitcell_array
Xport_data0 rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 dout0_32 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 din0_32 sel0_0 sel0_1 sel0_2 sel0_3 s_en0 p_en_bar0 w_en0 bank_wmask0_0 bank_wmask0_1 bank_wmask0_2 bank_wmask0_3 bank_spare_wen0_0 vdd gnd port_data
Xport_address0 addr0_2 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 addr0_8 addr0_9 wl_en0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 wl_0_128 rbl_wl0 vdd gnd port_address
Xcol_address_decoder0 addr0_0 addr0_1 sel0_0 sel0_1 sel0_2 sel0_3 vdd gnd hierarchical_predecode2x4_0
.ENDS bank
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* SPICE3 file created from sky130_fd_bd_sram__openram_dff.ext - technology: EFS8A

.subckt sky130_fd_bd_sram__openram_dff D Q CLK VDD GND
X1000 a_511_725# a_n8_115# VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1001 a_353_115# CLK a_11_624# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1002 a_353_725# a_203_89# a_11_624# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1003 a_11_624# a_203_89# a_161_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1004 a_11_624# CLK a_161_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1005 GND Q a_703_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1006 VDD Q a_703_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1007 a_203_89# CLK GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1008 a_203_89# CLK VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1009 a_161_115# D GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1010 a_161_725# D VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1011 GND a_11_624# a_n8_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1012 a_703_115# a_203_89# ON GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1013 VDD a_11_624# a_n8_115# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1014 a_703_725# CLK ON VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1015 Q ON VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1016 Q ON GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1017 ON a_203_89# a_511_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1018 ON CLK a_511_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1019 GND a_n8_115# a_353_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1020 VDD a_n8_115# a_353_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1021 a_511_115# a_n8_115# GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
.ends

.SUBCKT row_addr_dff din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 clk vdd gnd
*.PININFO din_0:I din_1:I din_2:I din_3:I din_4:I din_5:I din_6:I din_7:I dout_0:O dout_1:O dout_2:O dout_3:O dout_4:O dout_5:O dout_6:O dout_7:O clk:I vdd:B gnd:B
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 8 cols: 1
Xdff_r0_c0 din_0 dout_0 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r1_c0 din_1 dout_1 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r2_c0 din_2 dout_2 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r3_c0 din_3 dout_3 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r4_c0 din_4 dout_4 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r5_c0 din_5 dout_5 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r6_c0 din_6 dout_6 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r7_c0 din_7 dout_7 CLK VDD GND sky130_fd_bd_sram__openram_dff
.ENDS row_addr_dff

.SUBCKT col_addr_dff din_0 din_1 dout_0 dout_1 clk vdd gnd
*.PININFO din_0:I din_1:I dout_0:O dout_1:O clk:I vdd:B gnd:B
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 2
Xdff_r0_c0 din_0 dout_0 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c1 din_1 dout_1 CLK VDD GND sky130_fd_bd_sram__openram_dff
.ENDS col_addr_dff

.SUBCKT data_dff din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 din_32 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 dout_32 clk vdd gnd
*.PININFO din_0:I din_1:I din_2:I din_3:I din_4:I din_5:I din_6:I din_7:I din_8:I din_9:I din_10:I din_11:I din_12:I din_13:I din_14:I din_15:I din_16:I din_17:I din_18:I din_19:I din_20:I din_21:I din_22:I din_23:I din_24:I din_25:I din_26:I din_27:I din_28:I din_29:I din_30:I din_31:I din_32:I dout_0:O dout_1:O dout_2:O dout_3:O dout_4:O dout_5:O dout_6:O dout_7:O dout_8:O dout_9:O dout_10:O dout_11:O dout_12:O dout_13:O dout_14:O dout_15:O dout_16:O dout_17:O dout_18:O dout_19:O dout_20:O dout_21:O dout_22:O dout_23:O dout_24:O dout_25:O dout_26:O dout_27:O dout_28:O dout_29:O dout_30:O dout_31:O dout_32:O clk:I vdd:B gnd:B
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : din_32 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* OUTPUT: dout_32 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 33
Xdff_r0_c0 din_0 dout_0 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c1 din_1 dout_1 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c2 din_2 dout_2 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c3 din_3 dout_3 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c4 din_4 dout_4 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c5 din_5 dout_5 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c6 din_6 dout_6 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c7 din_7 dout_7 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c8 din_8 dout_8 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c9 din_9 dout_9 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c10 din_10 dout_10 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c11 din_11 dout_11 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c12 din_12 dout_12 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c13 din_13 dout_13 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c14 din_14 dout_14 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c15 din_15 dout_15 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c16 din_16 dout_16 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c17 din_17 dout_17 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c18 din_18 dout_18 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c19 din_19 dout_19 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c20 din_20 dout_20 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c21 din_21 dout_21 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c22 din_22 dout_22 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c23 din_23 dout_23 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c24 din_24 dout_24 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c25 din_25 dout_25 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c26 din_26 dout_26 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c27 din_27 dout_27 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c28 din_28 dout_28 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c29 din_29 dout_29 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c30 din_30 dout_30 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c31 din_31 dout_31 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c32 din_32 dout_32 CLK VDD GND sky130_fd_bd_sram__openram_dff
.ENDS data_dff

.SUBCKT wmask_dff din_0 din_1 din_2 din_3 dout_0 dout_1 dout_2 dout_3 clk vdd gnd
*.PININFO din_0:I din_1:I din_2:I din_3:I dout_0:O dout_1:O dout_2:O dout_3:O clk:I vdd:B gnd:B
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 4
Xdff_r0_c0 din_0 dout_0 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c1 din_1 dout_1 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c2 din_2 dout_2 CLK VDD GND sky130_fd_bd_sram__openram_dff
Xdff_r0_c3 din_3 dout_3 CLK VDD GND sky130_fd_bd_sram__openram_dff
.ENDS wmask_dff

.SUBCKT spare_wen_dff din_0 dout_0 clk vdd gnd
*.PININFO din_0:I dout_0:O clk:I vdd:B gnd:B
* INPUT : din_0 
* OUTPUT: dout_0 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 1
Xdff_r0_c0 din_0 dout_0 CLK VDD GND sky130_fd_bd_sram__openram_dff
.ENDS spare_wen_dff

.SUBCKT pinv_2 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=2 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pinv_2

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=3 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=3 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u

.SUBCKT pinv_3 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=3 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=3 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
.ENDS pinv_3

.SUBCKT dff_buf_0 D Q Qb clk vdd gnd
*.PININFO D:I Q:O Qb:O clk:I vdd:B gnd:B
* INPUT : D 
* OUTPUT: Q 
* OUTPUT: Qb 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_buf_dff D qint clk vdd gnd sky130_fd_bd_sram__openram_dff
Xdff_buf_inv1 qint Qb vdd gnd pinv_2
Xdff_buf_inv2 Qb Q vdd gnd pinv_3
.ENDS dff_buf_0

.SUBCKT dff_buf_array din_0 din_1 dout_0 dout_bar_0 dout_1 dout_bar_1 clk vdd gnd
*.PININFO din_0:I din_1:I dout_0:O dout_bar_0:O dout_1:O dout_bar_1:O clk:I vdd:B gnd:B
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_bar_0 
* OUTPUT: dout_1 
* OUTPUT: dout_bar_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_r0_c0 din_0 dout_0 dout_bar_0 clk vdd gnd dff_buf_0
Xdff_r1_c0 din_1 dout_1 dout_bar_1 clk vdd gnd dff_buf_0
.ENDS dff_buf_array

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=7 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=7 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_4 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=7 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=7 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
.ENDS pinv_4

.SUBCKT pdriver_1 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [12]
Xbuf_inv1 A Z vdd gnd pinv_4
.ENDS pdriver_1

.SUBCKT pand2_1 A B Z vdd gnd
*.PININFO A:I B:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand2_nand A B zb_int vdd gnd pnand2_0
Xpand2_inv zb_int Z vdd gnd pdriver_1
.ENDS pand2_1

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=18 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=18 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_5 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=18 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=18 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_5

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=70 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=70 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_6 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=70 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=70 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_6

.SUBCKT pbuf A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xbuf_inv1 A zb_int vdd gnd pinv_5
Xbuf_inv2 zb_int Z vdd gnd pinv_6
.ENDS pbuf

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=2 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_7 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=2 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u
.ENDS pinv_7

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=5 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=5 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_8 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=5 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=5 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_8

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=15 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=15 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_9 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=15 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=15 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_9

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=43 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=43 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_10 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=43 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=43 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_10

.SUBCKT pdriver_2 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 3, 9, 26, 78]
Xbuf_inv1 A Zb1_int vdd gnd pinv_0
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_0
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_7
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_8
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_9
Xbuf_inv6 Zb5_int Z vdd gnd pinv_10
.ENDS pdriver_2

.SUBCKT pinv_11 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=2 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pinv_11

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=3 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=3 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_12 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=3 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=3 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_12

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=8 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=8 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_13 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=8 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=8 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_13

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=24 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=24 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_14 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=24 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=24 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_14

.SUBCKT pdriver_3 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 2, 5, 14, 43]
Xbuf_inv1 A Zb1_int vdd gnd pinv_0
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_0
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_11
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_12
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_13
Xbuf_inv6 Zb5_int Z vdd gnd pinv_14
.ENDS pdriver_3

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

.SUBCKT pnand3 A B C Z vdd gnd
*.PININFO A:I B:I C:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpnand3_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand3_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand3_pmos3 Z C vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand3_nmos1 Z C net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand3_nmos2 net1 B net2 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand3_nmos3 net2 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pnand3

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=22 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=22 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_15 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=22 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=22 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_15

.SUBCKT pdriver_4 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [40]
Xbuf_inv1 A Z vdd gnd pinv_15
.ENDS pdriver_4

.SUBCKT pand3 A B C Z vdd gnd
*.PININFO A:I B:I C:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand A B C zb_int vdd gnd pnand3
Xpand3_inv zb_int Z vdd gnd pdriver_4
.ENDS pand3

.SUBCKT pinv_16 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=18 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=18 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_16

.SUBCKT pdriver_5 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [33]
Xbuf_inv1 A Z vdd gnd pinv_16
.ENDS pdriver_5

.SUBCKT pand3_0 A B C Z vdd gnd
*.PININFO A:I B:I C:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand A B C zb_int vdd gnd pnand3
Xpand3_inv zb_int Z vdd gnd pdriver_5
.ENDS pand3_0

.SUBCKT pnand2_1 A B Z vdd gnd
*.PININFO A:I B:I Z:O vdd:B gnd:B
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpnand2_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_nmos1 Z B net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand2_nmos2 net1 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pnand2_1

.SUBCKT pinv_17 A Z vdd gnd
*.PININFO A:I Z:O vdd:B gnd:B
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS pinv_17

.SUBCKT delay_chain in out vdd gnd
*.PININFO in:I out:O vdd:B gnd:B
* INPUT : in 
* OUTPUT: out 
* POWER : vdd 
* GROUND: gnd 
* fanouts: [4, 4, 4, 4, 4, 4, 4, 4, 4]
Xdinv0 in dout_1 vdd gnd pinv_17
Xdload_0_0 dout_1 n_0_0 vdd gnd pinv_17
Xdload_0_1 dout_1 n_0_1 vdd gnd pinv_17
Xdload_0_2 dout_1 n_0_2 vdd gnd pinv_17
Xdload_0_3 dout_1 n_0_3 vdd gnd pinv_17
Xdinv1 dout_1 dout_2 vdd gnd pinv_17
Xdload_1_0 dout_2 n_1_0 vdd gnd pinv_17
Xdload_1_1 dout_2 n_1_1 vdd gnd pinv_17
Xdload_1_2 dout_2 n_1_2 vdd gnd pinv_17
Xdload_1_3 dout_2 n_1_3 vdd gnd pinv_17
Xdinv2 dout_2 dout_3 vdd gnd pinv_17
Xdload_2_0 dout_3 n_2_0 vdd gnd pinv_17
Xdload_2_1 dout_3 n_2_1 vdd gnd pinv_17
Xdload_2_2 dout_3 n_2_2 vdd gnd pinv_17
Xdload_2_3 dout_3 n_2_3 vdd gnd pinv_17
Xdinv3 dout_3 dout_4 vdd gnd pinv_17
Xdload_3_0 dout_4 n_3_0 vdd gnd pinv_17
Xdload_3_1 dout_4 n_3_1 vdd gnd pinv_17
Xdload_3_2 dout_4 n_3_2 vdd gnd pinv_17
Xdload_3_3 dout_4 n_3_3 vdd gnd pinv_17
Xdinv4 dout_4 dout_5 vdd gnd pinv_17
Xdload_4_0 dout_5 n_4_0 vdd gnd pinv_17
Xdload_4_1 dout_5 n_4_1 vdd gnd pinv_17
Xdload_4_2 dout_5 n_4_2 vdd gnd pinv_17
Xdload_4_3 dout_5 n_4_3 vdd gnd pinv_17
Xdinv5 dout_5 dout_6 vdd gnd pinv_17
Xdload_5_0 dout_6 n_5_0 vdd gnd pinv_17
Xdload_5_1 dout_6 n_5_1 vdd gnd pinv_17
Xdload_5_2 dout_6 n_5_2 vdd gnd pinv_17
Xdload_5_3 dout_6 n_5_3 vdd gnd pinv_17
Xdinv6 dout_6 dout_7 vdd gnd pinv_17
Xdload_6_0 dout_7 n_6_0 vdd gnd pinv_17
Xdload_6_1 dout_7 n_6_1 vdd gnd pinv_17
Xdload_6_2 dout_7 n_6_2 vdd gnd pinv_17
Xdload_6_3 dout_7 n_6_3 vdd gnd pinv_17
Xdinv7 dout_7 dout_8 vdd gnd pinv_17
Xdload_7_0 dout_8 n_7_0 vdd gnd pinv_17
Xdload_7_1 dout_8 n_7_1 vdd gnd pinv_17
Xdload_7_2 dout_8 n_7_2 vdd gnd pinv_17
Xdload_7_3 dout_8 n_7_3 vdd gnd pinv_17
Xdinv8 dout_8 out vdd gnd pinv_17
Xdload_8_0 out n_8_0 vdd gnd pinv_17
Xdload_8_1 out n_8_1 vdd gnd pinv_17
Xdload_8_2 out n_8_2 vdd gnd pinv_17
Xdload_8_3 out n_8_3 vdd gnd pinv_17
.ENDS delay_chain

.SUBCKT control_logic_rw csb web clk rbl_bl s_en w_en p_en_bar wl_en clk_buf vdd gnd
*.PININFO csb:I web:I clk:I rbl_bl:I s_en:O w_en:O p_en_bar:O wl_en:O clk_buf:O vdd:B gnd:B
* INPUT : csb 
* INPUT : web 
* INPUT : clk 
* INPUT : rbl_bl 
* OUTPUT: s_en 
* OUTPUT: w_en 
* OUTPUT: p_en_bar 
* OUTPUT: wl_en 
* OUTPUT: clk_buf 
* POWER : vdd 
* GROUND: gnd 
* word_size 32
Xctrl_dffs csb web cs_bar cs we_bar we clk_buf vdd gnd dff_buf_array
Xclkbuf clk clk_buf vdd gnd pdriver_2
Xinv_clk_bar clk_buf clk_bar vdd gnd pinv_1
Xand2_gated_clk_bar clk_bar cs gated_clk_bar vdd gnd pand2_1
Xand2_gated_clk_buf clk_buf cs gated_clk_buf vdd gnd pand2_1
Xbuf_wl_en gated_clk_bar wl_en vdd gnd pdriver_3
Xrbl_bl_delay_inv rbl_bl_delay rbl_bl_delay_bar vdd gnd pinv_1
Xw_en_and we rbl_bl_delay_bar gated_clk_bar w_en vdd gnd pand3
Xbuf_s_en_and rbl_bl_delay gated_clk_bar we_bar s_en vdd gnd pand3_0
Xdelay_chain rbl_bl rbl_bl_delay vdd gnd delay_chain
Xnand_p_en_bar gated_clk_buf rbl_bl_delay p_en_bar_unbuf vdd gnd pnand2_1
Xbuf_p_en_bar p_en_bar_unbuf p_en_bar vdd gnd pdriver_3
.ENDS control_logic_rw

.SUBCKT sky130_sram_2kbyte_1rw_32x512_8 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] din0[32] addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] addr0[9] csb0 web0 clk0 wmask0[0] wmask0[1] wmask0[2] wmask0[3] spare_wen0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] dout0[32] vccd1 vssd1
*.PININFO din0[0]:I din0[1]:I din0[2]:I din0[3]:I din0[4]:I din0[5]:I din0[6]:I din0[7]:I din0[8]:I din0[9]:I din0[10]:I din0[11]:I din0[12]:I din0[13]:I din0[14]:I din0[15]:I din0[16]:I din0[17]:I din0[18]:I din0[19]:I din0[20]:I din0[21]:I din0[22]:I din0[23]:I din0[24]:I din0[25]:I din0[26]:I din0[27]:I din0[28]:I din0[29]:I din0[30]:I din0[31]:I din0[32]:I addr0[0]:I addr0[1]:I addr0[2]:I addr0[3]:I addr0[4]:I addr0[5]:I addr0[6]:I addr0[7]:I addr0[8]:I addr0[9]:I csb0:I web0:I clk0:I wmask0[0]:I wmask0[1]:I wmask0[2]:I wmask0[3]:I spare_wen0:I dout0[0]:O dout0[1]:O dout0[2]:O dout0[3]:O dout0[4]:O dout0[5]:O dout0[6]:O dout0[7]:O dout0[8]:O dout0[9]:O dout0[10]:O dout0[11]:O dout0[12]:O dout0[13]:O dout0[14]:O dout0[15]:O dout0[16]:O dout0[17]:O dout0[18]:O dout0[19]:O dout0[20]:O dout0[21]:O dout0[22]:O dout0[23]:O dout0[24]:O dout0[25]:O dout0[26]:O dout0[27]:O dout0[28]:O dout0[29]:O dout0[30]:O dout0[31]:O dout0[32]:O vccd1:B vssd1:B
* INPUT : din0[0] 
* INPUT : din0[1] 
* INPUT : din0[2] 
* INPUT : din0[3] 
* INPUT : din0[4] 
* INPUT : din0[5] 
* INPUT : din0[6] 
* INPUT : din0[7] 
* INPUT : din0[8] 
* INPUT : din0[9] 
* INPUT : din0[10] 
* INPUT : din0[11] 
* INPUT : din0[12] 
* INPUT : din0[13] 
* INPUT : din0[14] 
* INPUT : din0[15] 
* INPUT : din0[16] 
* INPUT : din0[17] 
* INPUT : din0[18] 
* INPUT : din0[19] 
* INPUT : din0[20] 
* INPUT : din0[21] 
* INPUT : din0[22] 
* INPUT : din0[23] 
* INPUT : din0[24] 
* INPUT : din0[25] 
* INPUT : din0[26] 
* INPUT : din0[27] 
* INPUT : din0[28] 
* INPUT : din0[29] 
* INPUT : din0[30] 
* INPUT : din0[31] 
* INPUT : din0[32] 
* INPUT : addr0[0] 
* INPUT : addr0[1] 
* INPUT : addr0[2] 
* INPUT : addr0[3] 
* INPUT : addr0[4] 
* INPUT : addr0[5] 
* INPUT : addr0[6] 
* INPUT : addr0[7] 
* INPUT : addr0[8] 
* INPUT : addr0[9] 
* INPUT : csb0 
* INPUT : web0 
* INPUT : clk0 
* INPUT : wmask0[0] 
* INPUT : wmask0[1] 
* INPUT : wmask0[2] 
* INPUT : wmask0[3] 
* INPUT : spare_wen0 
* OUTPUT: dout0[0] 
* OUTPUT: dout0[1] 
* OUTPUT: dout0[2] 
* OUTPUT: dout0[3] 
* OUTPUT: dout0[4] 
* OUTPUT: dout0[5] 
* OUTPUT: dout0[6] 
* OUTPUT: dout0[7] 
* OUTPUT: dout0[8] 
* OUTPUT: dout0[9] 
* OUTPUT: dout0[10] 
* OUTPUT: dout0[11] 
* OUTPUT: dout0[12] 
* OUTPUT: dout0[13] 
* OUTPUT: dout0[14] 
* OUTPUT: dout0[15] 
* OUTPUT: dout0[16] 
* OUTPUT: dout0[17] 
* OUTPUT: dout0[18] 
* OUTPUT: dout0[19] 
* OUTPUT: dout0[20] 
* OUTPUT: dout0[21] 
* OUTPUT: dout0[22] 
* OUTPUT: dout0[23] 
* OUTPUT: dout0[24] 
* OUTPUT: dout0[25] 
* OUTPUT: dout0[26] 
* OUTPUT: dout0[27] 
* OUTPUT: dout0[28] 
* OUTPUT: dout0[29] 
* OUTPUT: dout0[30] 
* OUTPUT: dout0[31] 
* OUTPUT: dout0[32] 
* POWER : vccd1 
* GROUND: vssd1 
Xbank0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] dout0[32] rbl_bl0 bank_din0_0 bank_din0_1 bank_din0_2 bank_din0_3 bank_din0_4 bank_din0_5 bank_din0_6 bank_din0_7 bank_din0_8 bank_din0_9 bank_din0_10 bank_din0_11 bank_din0_12 bank_din0_13 bank_din0_14 bank_din0_15 bank_din0_16 bank_din0_17 bank_din0_18 bank_din0_19 bank_din0_20 bank_din0_21 bank_din0_22 bank_din0_23 bank_din0_24 bank_din0_25 bank_din0_26 bank_din0_27 bank_din0_28 bank_din0_29 bank_din0_30 bank_din0_31 bank_din0_32 a0_0 a0_1 a0_2 a0_3 a0_4 a0_5 a0_6 a0_7 a0_8 a0_9 s_en0 p_en_bar0 w_en0 bank_wmask0_0 bank_wmask0_1 bank_wmask0_2 bank_wmask0_3 bank_spare_wen0_0 wl_en0 vccd1 vssd1 bank
Xcontrol0 csb0 web0 clk0 rbl_bl0 s_en0 w_en0 p_en_bar0 wl_en0 clk_buf0 vccd1 vssd1 control_logic_rw
Xrow_address0 addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] addr0[9] a0_2 a0_3 a0_4 a0_5 a0_6 a0_7 a0_8 a0_9 clk_buf0 vccd1 vssd1 row_addr_dff
Xcol_address0 addr0[0] addr0[1] a0_0 a0_1 clk_buf0 vccd1 vssd1 col_addr_dff
Xwmask_dff0 wmask0[0] wmask0[1] wmask0[2] wmask0[3] bank_wmask0_0 bank_wmask0_1 bank_wmask0_2 bank_wmask0_3 clk_buf0 vccd1 vssd1 wmask_dff
Xdata_dff0 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] din0[32] bank_din0_0 bank_din0_1 bank_din0_2 bank_din0_3 bank_din0_4 bank_din0_5 bank_din0_6 bank_din0_7 bank_din0_8 bank_din0_9 bank_din0_10 bank_din0_11 bank_din0_12 bank_din0_13 bank_din0_14 bank_din0_15 bank_din0_16 bank_din0_17 bank_din0_18 bank_din0_19 bank_din0_20 bank_din0_21 bank_din0_22 bank_din0_23 bank_din0_24 bank_din0_25 bank_din0_26 bank_din0_27 bank_din0_28 bank_din0_29 bank_din0_30 bank_din0_31 bank_din0_32 clk_buf0 vccd1 vssd1 data_dff
Xspare_wen_dff0 spare_wen0[0] bank_spare_wen0_0 clk_buf0 vccd1 vssd1 spare_wen_dff
.ENDS sky130_sram_2kbyte_1rw_32x512_8
