VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_1kbyte_1rw1r_8x1024_8
   CLASS BLOCK ;
   SIZE 437.62 BY 432.18 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.24 0.0 80.62 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  86.36 0.0 86.74 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.8 0.0 92.18 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  97.24 0.0 97.62 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  103.36 0.0 103.74 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.8 0.0 109.18 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  115.6 0.0 115.98 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  120.36 0.0 120.74 0.38 ;
      END
   END din0[7]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  56.44 0.0 56.82 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  63.24 0.0 63.62 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  68.68 0.0 69.06 0.38 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 136.0 0.38 136.38 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 144.16 0.38 144.54 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 150.96 0.38 151.34 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 159.12 0.38 159.5 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 164.56 0.38 164.94 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 172.72 0.38 173.1 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 178.16 0.38 178.54 ;
      END
   END addr0[9]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  375.36 431.8 375.74 432.18 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  369.92 431.8 370.3 432.18 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  364.48 431.8 364.86 432.18 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  437.24 91.8 437.62 92.18 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  437.24 82.96 437.62 83.34 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  437.24 77.52 437.62 77.9 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  437.24 68.68 437.62 69.06 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  437.24 63.24 437.62 63.62 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  437.24 55.08 437.62 55.46 ;
      END
   END addr1[8]
   PIN addr1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  437.24 48.28 437.62 48.66 ;
      END
   END addr1[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 36.04 0.38 36.42 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  437.24 390.32 437.62 390.7 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 44.2 0.38 44.58 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 36.72 0.38 37.1 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  437.24 389.64 437.62 390.02 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  74.12 0.0 74.5 0.38 ;
      END
   END wmask0[0]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  118.32 0.0 118.7 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  144.16 0.0 144.54 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  169.32 0.0 169.7 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  194.48 0.0 194.86 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  219.64 0.0 220.02 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  244.12 0.0 244.5 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.28 0.0 269.66 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  294.44 0.0 294.82 0.38 ;
      END
   END dout0[7]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  119.68 431.8 120.06 432.18 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  144.84 431.8 145.22 432.18 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  170.0 431.8 170.38 432.18 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  195.16 431.8 195.54 432.18 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  219.64 431.8 220.02 432.18 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  244.12 431.8 244.5 432.18 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.96 431.8 270.34 432.18 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  295.12 431.8 295.5 432.18 ;
      END
   END dout1[7]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  1.36 0.0 2.42 431.5 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.06 431.5 ;
      END
   END gnd
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 437.0 431.56 ;
   LAYER  met2 ;
      RECT  0.62 0.62 437.0 431.56 ;
   LAYER  met3 ;
      RECT  0.68 135.7 437.0 136.68 ;
      RECT  0.62 136.68 0.68 143.86 ;
      RECT  0.62 144.84 0.68 150.66 ;
      RECT  0.62 151.64 0.68 158.82 ;
      RECT  0.62 159.8 0.68 164.26 ;
      RECT  0.62 165.24 0.68 172.42 ;
      RECT  0.62 173.4 0.68 177.86 ;
      RECT  0.62 178.84 0.68 431.56 ;
      RECT  0.68 0.62 436.94 91.5 ;
      RECT  0.68 91.5 436.94 92.48 ;
      RECT  0.68 92.48 436.94 135.7 ;
      RECT  436.94 92.48 437.0 135.7 ;
      RECT  436.94 83.64 437.0 91.5 ;
      RECT  436.94 78.2 437.0 82.66 ;
      RECT  436.94 69.36 437.0 77.22 ;
      RECT  436.94 63.92 437.0 68.38 ;
      RECT  436.94 55.76 437.0 62.94 ;
      RECT  436.94 0.62 437.0 47.98 ;
      RECT  436.94 48.96 437.0 54.78 ;
      RECT  0.62 0.62 0.68 35.74 ;
      RECT  0.68 136.68 436.94 390.02 ;
      RECT  0.68 390.02 436.94 391.0 ;
      RECT  0.68 391.0 436.94 431.56 ;
      RECT  436.94 391.0 437.0 431.56 ;
      RECT  0.62 44.88 0.68 135.7 ;
      RECT  0.62 37.4 0.68 43.9 ;
      RECT  436.94 136.68 437.0 389.34 ;
   LAYER  met4 ;
      RECT  79.94 0.68 80.92 431.56 ;
      RECT  80.92 0.62 86.06 0.68 ;
      RECT  87.04 0.62 91.5 0.68 ;
      RECT  92.48 0.62 96.94 0.68 ;
      RECT  97.92 0.62 103.06 0.68 ;
      RECT  104.04 0.62 108.5 0.68 ;
      RECT  109.48 0.62 115.3 0.68 ;
      RECT  57.12 0.62 62.94 0.68 ;
      RECT  63.92 0.62 68.38 0.68 ;
      RECT  80.92 0.68 375.06 431.5 ;
      RECT  375.06 0.68 376.04 431.5 ;
      RECT  376.04 0.68 437.0 431.5 ;
      RECT  376.04 431.5 437.0 431.56 ;
      RECT  370.6 431.5 375.06 431.56 ;
      RECT  365.16 431.5 369.62 431.56 ;
      RECT  69.36 0.62 73.82 0.68 ;
      RECT  74.8 0.62 79.94 0.68 ;
      RECT  116.28 0.62 118.02 0.68 ;
      RECT  119.0 0.62 120.06 0.68 ;
      RECT  121.04 0.62 143.86 0.68 ;
      RECT  144.84 0.62 169.02 0.68 ;
      RECT  170.0 0.62 194.18 0.68 ;
      RECT  195.16 0.62 219.34 0.68 ;
      RECT  220.32 0.62 243.82 0.68 ;
      RECT  244.8 0.62 268.98 0.68 ;
      RECT  269.96 0.62 294.14 0.68 ;
      RECT  295.12 0.62 437.0 0.68 ;
      RECT  80.92 431.5 119.38 431.56 ;
      RECT  120.36 431.5 144.54 431.56 ;
      RECT  145.52 431.5 169.7 431.56 ;
      RECT  170.68 431.5 194.86 431.56 ;
      RECT  195.84 431.5 219.34 431.56 ;
      RECT  220.32 431.5 243.82 431.56 ;
      RECT  244.8 431.5 269.66 431.56 ;
      RECT  270.64 431.5 294.82 431.56 ;
      RECT  295.8 431.5 364.18 431.56 ;
      RECT  2.72 0.68 79.94 431.56 ;
      RECT  2.72 0.62 56.14 0.68 ;
   END
END    sky130_sram_1kbyte_1rw1r_8x1024_8
END    LIBRARY
